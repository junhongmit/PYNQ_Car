----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:05:12 03/26/2014 
-- Design Name: 
-- Module Name:    LineBuffer - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LineBuffer_vhdl is
port(
clock:		in 		std_logic;
clken,aclr: in 		std_logic;
shiftin:		in 		std_logic_vector(7 downto 0);
shiftout:	out 		std_logic_vector(7 downto 0);
taps:			out 		std_logic_vector(23 downto 0)
);
end LineBuffer_vhdl;

architecture Behavioral of LineBuffer_vhdl is


subtype word is std_logic_vector(7 downto 0);
type memory is array(0 to 1279)of word;
signal LineBuffer0:memory;
signal LineBuffer1:memory;
signal LineBuffer2:memory;
signal taps_signal :	std_logic_vector(23 downto 0);
begin

process(clock,aclr,clken)
begin

 if(clken = '1')then
   if rising_edge(clock)then
         if(aclr = '1')then
			LineBuffer0(0) <= "00000000";
			LineBuffer0(1) <= "00000000";
			LineBuffer0(2) <= "00000000";
			LineBuffer0(3) <= "00000000";
			LineBuffer0(4) <= "00000000";
			LineBuffer0(5) <= "00000000";
			LineBuffer0(6) <= "00000000";
			LineBuffer0(7) <= "00000000";
			LineBuffer0(8) <= "00000000";
			LineBuffer0(9) <= "00000000";	
			LineBuffer0(10) <= "00000000";
			LineBuffer0(11) <= "00000000";
			LineBuffer0(12) <= "00000000";
			LineBuffer0(13) <= "00000000";
			LineBuffer0(14) <= "00000000";
			LineBuffer0(15) <= "00000000";
			LineBuffer0(16) <= "00000000";
			LineBuffer0(17) <= "00000000";
			LineBuffer0(18) <= "00000000";
			LineBuffer0(19) <= "00000000";	
			LineBuffer0(20) <= "00000000";
			LineBuffer0(21) <= "00000000";
			LineBuffer0(22) <= "00000000";
			LineBuffer0(23) <= "00000000";
			LineBuffer0(24) <= "00000000";
			LineBuffer0(25) <= "00000000";
			LineBuffer0(26) <= "00000000";
			LineBuffer0(27) <= "00000000";
			LineBuffer0(28) <= "00000000";
			LineBuffer0(29) <= "00000000";	
			LineBuffer0(30) <= "00000000";
			LineBuffer0(31) <= "00000000";
			LineBuffer0(32) <= "00000000";
			LineBuffer0(33) <= "00000000";
			LineBuffer0(34) <= "00000000";
			LineBuffer0(35) <= "00000000";
			LineBuffer0(36) <= "00000000";
			LineBuffer0(37) <= "00000000";
			LineBuffer0(38) <= "00000000";
			LineBuffer0(39) <= "00000000";	
			LineBuffer0(40) <= "00000000";
			LineBuffer0(41) <= "00000000";
			LineBuffer0(42) <= "00000000";
			LineBuffer0(43) <= "00000000";
			LineBuffer0(44) <= "00000000";
			LineBuffer0(45) <= "00000000";
			LineBuffer0(46) <= "00000000";
			LineBuffer0(47) <= "00000000";
			LineBuffer0(48) <= "00000000";
			LineBuffer0(49) <= "00000000";	
			LineBuffer0(50) <= "00000000";
			LineBuffer0(51) <= "00000000";
			LineBuffer0(52) <= "00000000";
			LineBuffer0(53) <= "00000000";
			LineBuffer0(54) <= "00000000";
			LineBuffer0(55) <= "00000000";
			LineBuffer0(56) <= "00000000";
			LineBuffer0(57) <= "00000000";
			LineBuffer0(58) <= "00000000";
			LineBuffer0(59) <= "00000000";	
			LineBuffer0(60) <= "00000000";
			LineBuffer0(61) <= "00000000";
			LineBuffer0(62) <= "00000000";
			LineBuffer0(63) <= "00000000";
			LineBuffer0(64) <= "00000000";
			LineBuffer0(65) <= "00000000";
			LineBuffer0(66) <= "00000000";
			LineBuffer0(67) <= "00000000";
			LineBuffer0(68) <= "00000000";
			LineBuffer0(69) <= "00000000";	
			LineBuffer0(70) <= "00000000";
			LineBuffer0(71) <= "00000000";
			LineBuffer0(72) <= "00000000";
			LineBuffer0(73) <= "00000000";
			LineBuffer0(74) <= "00000000";
			LineBuffer0(75) <= "00000000";
			LineBuffer0(76) <= "00000000";
			LineBuffer0(77) <= "00000000";
			LineBuffer0(78) <= "00000000";
			LineBuffer0(79) <= "00000000";	
			LineBuffer0(80) <= "00000000";
			LineBuffer0(81) <= "00000000";
			LineBuffer0(82) <= "00000000";
			LineBuffer0(83) <= "00000000";
			LineBuffer0(84) <= "00000000";
			LineBuffer0(85) <= "00000000";
			LineBuffer0(86) <= "00000000";
			LineBuffer0(87) <= "00000000";
			LineBuffer0(88) <= "00000000";
			LineBuffer0(89) <= "00000000";	
			LineBuffer0(90) <= "00000000";
			LineBuffer0(91) <= "00000000";
			LineBuffer0(92) <= "00000000";
			LineBuffer0(93) <= "00000000";
			LineBuffer0(94) <= "00000000";
			LineBuffer0(95) <= "00000000";
			LineBuffer0(96) <= "00000000";
			LineBuffer0(97) <= "00000000";
			LineBuffer0(98) <= "00000000";
			LineBuffer0(99) <= "00000000";	
			LineBuffer0(100) <= "00000000";
			LineBuffer0(101) <= "00000000";
			LineBuffer0(102) <= "00000000";
			LineBuffer0(103) <= "00000000";
			LineBuffer0(104) <= "00000000";
			LineBuffer0(105) <= "00000000";
			LineBuffer0(106) <= "00000000";
			LineBuffer0(107) <= "00000000";
			LineBuffer0(108) <= "00000000";
			LineBuffer0(109) <= "00000000";	
			LineBuffer0(110) <= "00000000";
			LineBuffer0(111) <= "00000000";
			LineBuffer0(112) <= "00000000";
			LineBuffer0(113) <= "00000000";
			LineBuffer0(114) <= "00000000";
			LineBuffer0(115) <= "00000000";
			LineBuffer0(116) <= "00000000";
			LineBuffer0(117) <= "00000000";
			LineBuffer0(118) <= "00000000";
			LineBuffer0(119) <= "00000000";	
			LineBuffer0(120) <= "00000000";
			LineBuffer0(121) <= "00000000";
			LineBuffer0(122) <= "00000000";
			LineBuffer0(123) <= "00000000";
			LineBuffer0(124) <= "00000000";
			LineBuffer0(125) <= "00000000";
			LineBuffer0(126) <= "00000000";
			LineBuffer0(127) <= "00000000";
			LineBuffer0(128) <= "00000000";
			LineBuffer0(129) <= "00000000";	
			LineBuffer0(130) <= "00000000";
			LineBuffer0(131) <= "00000000";
			LineBuffer0(132) <= "00000000";
			LineBuffer0(133) <= "00000000";
			LineBuffer0(134) <= "00000000";
			LineBuffer0(135) <= "00000000";
			LineBuffer0(136) <= "00000000";
			LineBuffer0(137) <= "00000000";
			LineBuffer0(138) <= "00000000";
			LineBuffer0(139) <= "00000000";	
			LineBuffer0(140) <= "00000000";
			LineBuffer0(141) <= "00000000";
			LineBuffer0(142) <= "00000000";
			LineBuffer0(143) <= "00000000";
			LineBuffer0(144) <= "00000000";
			LineBuffer0(145) <= "00000000";
			LineBuffer0(146) <= "00000000";
			LineBuffer0(147) <= "00000000";
			LineBuffer0(148) <= "00000000";
			LineBuffer0(149) <= "00000000";	
			LineBuffer0(150) <= "00000000";
			LineBuffer0(151) <= "00000000";
			LineBuffer0(152) <= "00000000";
			LineBuffer0(153) <= "00000000";
			LineBuffer0(154) <= "00000000";
			LineBuffer0(155) <= "00000000";
			LineBuffer0(156) <= "00000000";
			LineBuffer0(157) <= "00000000";
			LineBuffer0(158) <= "00000000";
			LineBuffer0(159) <= "00000000";	
			LineBuffer0(160) <= "00000000";
			LineBuffer0(161) <= "00000000";
			LineBuffer0(162) <= "00000000";
			LineBuffer0(163) <= "00000000";
			LineBuffer0(164) <= "00000000";
			LineBuffer0(165) <= "00000000";
			LineBuffer0(166) <= "00000000";
			LineBuffer0(167) <= "00000000";
			LineBuffer0(168) <= "00000000";
			LineBuffer0(169) <= "00000000";	
			LineBuffer0(170) <= "00000000";
			LineBuffer0(171) <= "00000000";
			LineBuffer0(172) <= "00000000";
			LineBuffer0(173) <= "00000000";
			LineBuffer0(174) <= "00000000";
			LineBuffer0(175) <= "00000000";
			LineBuffer0(176) <= "00000000";
			LineBuffer0(177) <= "00000000";
			LineBuffer0(178) <= "00000000";
			LineBuffer0(179) <= "00000000";	
			LineBuffer0(180) <= "00000000";
			LineBuffer0(181) <= "00000000";
			LineBuffer0(182) <= "00000000";
			LineBuffer0(183) <= "00000000";
			LineBuffer0(184) <= "00000000";
			LineBuffer0(185) <= "00000000";
			LineBuffer0(186) <= "00000000";
			LineBuffer0(187) <= "00000000";
			LineBuffer0(188) <= "00000000";
			LineBuffer0(189) <= "00000000";	
			LineBuffer0(190) <= "00000000";
			LineBuffer0(191) <= "00000000";
			LineBuffer0(192) <= "00000000";
			LineBuffer0(193) <= "00000000";
			LineBuffer0(194) <= "00000000";
			LineBuffer0(195) <= "00000000";
			LineBuffer0(196) <= "00000000";
			LineBuffer0(197) <= "00000000";
			LineBuffer0(198) <= "00000000";
			LineBuffer0(199) <= "00000000";
			LineBuffer0(200) <= "00000000";
			LineBuffer0(201) <= "00000000";
			LineBuffer0(202) <= "00000000";
			LineBuffer0(203) <= "00000000";
			LineBuffer0(204) <= "00000000";
			LineBuffer0(205) <= "00000000";
			LineBuffer0(206) <= "00000000";
			LineBuffer0(207) <= "00000000";
			LineBuffer0(208) <= "00000000";
			LineBuffer0(209) <= "00000000";	
			LineBuffer0(210) <= "00000000";
			LineBuffer0(211) <= "00000000";
			LineBuffer0(212) <= "00000000";
			LineBuffer0(213) <= "00000000";
			LineBuffer0(214) <= "00000000";
			LineBuffer0(215) <= "00000000";
			LineBuffer0(216) <= "00000000";
			LineBuffer0(217) <= "00000000";
			LineBuffer0(218) <= "00000000";
			LineBuffer0(219) <= "00000000";	
			LineBuffer0(220) <= "00000000";
			LineBuffer0(221) <= "00000000";
			LineBuffer0(222) <= "00000000";
			LineBuffer0(223) <= "00000000";
			LineBuffer0(224) <= "00000000";
			LineBuffer0(225) <= "00000000";
			LineBuffer0(226) <= "00000000";
			LineBuffer0(227) <= "00000000";
			LineBuffer0(228) <= "00000000";
			LineBuffer0(229) <= "00000000";	
			LineBuffer0(230) <= "00000000";
			LineBuffer0(231) <= "00000000";
			LineBuffer0(232) <= "00000000";
			LineBuffer0(233) <= "00000000";
			LineBuffer0(234) <= "00000000";
			LineBuffer0(235) <= "00000000";
			LineBuffer0(236) <= "00000000";
			LineBuffer0(237) <= "00000000";
			LineBuffer0(238) <= "00000000";
			LineBuffer0(239) <= "00000000";	
			LineBuffer0(240) <= "00000000";
			LineBuffer0(241) <= "00000000";
			LineBuffer0(242) <= "00000000";
			LineBuffer0(243) <= "00000000";
			LineBuffer0(244) <= "00000000";
			LineBuffer0(245) <= "00000000";
			LineBuffer0(246) <= "00000000";
			LineBuffer0(247) <= "00000000";
			LineBuffer0(248) <= "00000000";
			LineBuffer0(249) <= "00000000";	
			LineBuffer0(250) <= "00000000";
			LineBuffer0(251) <= "00000000";
			LineBuffer0(252) <= "00000000";
			LineBuffer0(253) <= "00000000";
			LineBuffer0(254) <= "00000000";
			LineBuffer0(255) <= "00000000";
			LineBuffer0(256) <= "00000000";
			LineBuffer0(257) <= "00000000";
			LineBuffer0(258) <= "00000000";
			LineBuffer0(259) <= "00000000";	
			LineBuffer0(260) <= "00000000";
			LineBuffer0(261) <= "00000000";
			LineBuffer0(262) <= "00000000";
			LineBuffer0(263) <= "00000000";
			LineBuffer0(264) <= "00000000";
			LineBuffer0(265) <= "00000000";
			LineBuffer0(266) <= "00000000";
			LineBuffer0(267) <= "00000000";
			LineBuffer0(268) <= "00000000";
			LineBuffer0(269) <= "00000000";	
			LineBuffer0(270) <= "00000000";
			LineBuffer0(271) <= "00000000";
			LineBuffer0(272) <= "00000000";
			LineBuffer0(273) <= "00000000";
			LineBuffer0(274) <= "00000000";
			LineBuffer0(275) <= "00000000";
			LineBuffer0(276) <= "00000000";
			LineBuffer0(277) <= "00000000";
			LineBuffer0(278) <= "00000000";
			LineBuffer0(279) <= "00000000";	
			LineBuffer0(280) <= "00000000";
			LineBuffer0(281) <= "00000000";
			LineBuffer0(282) <= "00000000";
			LineBuffer0(283) <= "00000000";
			LineBuffer0(284) <= "00000000";
			LineBuffer0(285) <= "00000000";
			LineBuffer0(286) <= "00000000";
			LineBuffer0(287) <= "00000000";
			LineBuffer0(288) <= "00000000";
			LineBuffer0(289) <= "00000000";	
			LineBuffer0(290) <= "00000000";
			LineBuffer0(291) <= "00000000";
			LineBuffer0(292) <= "00000000";
			LineBuffer0(293) <= "00000000";
			LineBuffer0(294) <= "00000000";
			LineBuffer0(295) <= "00000000";
			LineBuffer0(296) <= "00000000";
			LineBuffer0(297) <= "00000000";
			LineBuffer0(298) <= "00000000";
			LineBuffer0(299) <= "00000000";
			LineBuffer0(300) <= "00000000";
			LineBuffer0(301) <= "00000000";
			LineBuffer0(302) <= "00000000";
			LineBuffer0(303) <= "00000000";
			LineBuffer0(304) <= "00000000";
			LineBuffer0(305) <= "00000000";
			LineBuffer0(306) <= "00000000";
			LineBuffer0(307) <= "00000000";
			LineBuffer0(308) <= "00000000";
			LineBuffer0(309) <= "00000000";	
			LineBuffer0(310) <= "00000000";
			LineBuffer0(311) <= "00000000";
			LineBuffer0(312) <= "00000000";
			LineBuffer0(313) <= "00000000";
			LineBuffer0(314) <= "00000000";
			LineBuffer0(315) <= "00000000";
			LineBuffer0(316) <= "00000000";
			LineBuffer0(317) <= "00000000";
			LineBuffer0(318) <= "00000000";
			LineBuffer0(319) <= "00000000";	
			LineBuffer0(320) <= "00000000";
			LineBuffer0(321) <= "00000000";
			LineBuffer0(322) <= "00000000";
			LineBuffer0(323) <= "00000000";
			LineBuffer0(324) <= "00000000";
			LineBuffer0(325) <= "00000000";
			LineBuffer0(326) <= "00000000";
			LineBuffer0(327) <= "00000000";
			LineBuffer0(328) <= "00000000";
			LineBuffer0(329) <= "00000000";	
			LineBuffer0(330) <= "00000000";
			LineBuffer0(331) <= "00000000";
			LineBuffer0(332) <= "00000000";
			LineBuffer0(333) <= "00000000";
			LineBuffer0(334) <= "00000000";
			LineBuffer0(335) <= "00000000";
			LineBuffer0(336) <= "00000000";
			LineBuffer0(337) <= "00000000";
			LineBuffer0(338) <= "00000000";
			LineBuffer0(339) <= "00000000";	
			LineBuffer0(340) <= "00000000";
			LineBuffer0(341) <= "00000000";
			LineBuffer0(342) <= "00000000";
			LineBuffer0(343) <= "00000000";
			LineBuffer0(344) <= "00000000";
			LineBuffer0(345) <= "00000000";
			LineBuffer0(346) <= "00000000";
			LineBuffer0(347) <= "00000000";
			LineBuffer0(348) <= "00000000";
			LineBuffer0(349) <= "00000000";	
			LineBuffer0(350) <= "00000000";
			LineBuffer0(351) <= "00000000";
			LineBuffer0(352) <= "00000000";
			LineBuffer0(353) <= "00000000";
			LineBuffer0(354) <= "00000000";
			LineBuffer0(355) <= "00000000";
			LineBuffer0(356) <= "00000000";
			LineBuffer0(357) <= "00000000";
			LineBuffer0(358) <= "00000000";
			LineBuffer0(359) <= "00000000";	
			LineBuffer0(360) <= "00000000";
			LineBuffer0(361) <= "00000000";
			LineBuffer0(362) <= "00000000";
			LineBuffer0(363) <= "00000000";
			LineBuffer0(364) <= "00000000";
			LineBuffer0(365) <= "00000000";
			LineBuffer0(366) <= "00000000";
			LineBuffer0(367) <= "00000000";
			LineBuffer0(368) <= "00000000";
			LineBuffer0(369) <= "00000000";	
			LineBuffer0(370) <= "00000000";
			LineBuffer0(371) <= "00000000";
			LineBuffer0(372) <= "00000000";
			LineBuffer0(373) <= "00000000";
			LineBuffer0(374) <= "00000000";
			LineBuffer0(375) <= "00000000";
			LineBuffer0(376) <= "00000000";
			LineBuffer0(377) <= "00000000";
			LineBuffer0(378) <= "00000000";
			LineBuffer0(379) <= "00000000";	
			LineBuffer0(380) <= "00000000";
			LineBuffer0(381) <= "00000000";
			LineBuffer0(382) <= "00000000";
			LineBuffer0(383) <= "00000000";
			LineBuffer0(384) <= "00000000";
			LineBuffer0(385) <= "00000000";
			LineBuffer0(386) <= "00000000";
			LineBuffer0(387) <= "00000000";
			LineBuffer0(388) <= "00000000";
			LineBuffer0(389) <= "00000000";	
			LineBuffer0(390) <= "00000000";
			LineBuffer0(391) <= "00000000";
			LineBuffer0(392) <= "00000000";
			LineBuffer0(393) <= "00000000";
			LineBuffer0(394) <= "00000000";
			LineBuffer0(395) <= "00000000";
			LineBuffer0(396) <= "00000000";
			LineBuffer0(397) <= "00000000";
			LineBuffer0(398) <= "00000000";
			LineBuffer0(399) <= "00000000";
			LineBuffer0(400) <= "00000000";
			LineBuffer0(401) <= "00000000";
			LineBuffer0(402) <= "00000000";
			LineBuffer0(403) <= "00000000";
			LineBuffer0(404) <= "00000000";
			LineBuffer0(405) <= "00000000";
			LineBuffer0(406) <= "00000000";
			LineBuffer0(407) <= "00000000";
			LineBuffer0(408) <= "00000000";
			LineBuffer0(409) <= "00000000";	
			LineBuffer0(410) <= "00000000";
			LineBuffer0(411) <= "00000000";
			LineBuffer0(412) <= "00000000";
			LineBuffer0(413) <= "00000000";
			LineBuffer0(414) <= "00000000";
			LineBuffer0(415) <= "00000000";
			LineBuffer0(416) <= "00000000";
			LineBuffer0(417) <= "00000000";
			LineBuffer0(418) <= "00000000";
			LineBuffer0(419) <= "00000000";	
			LineBuffer0(420) <= "00000000";
			LineBuffer0(421) <= "00000000";
			LineBuffer0(422) <= "00000000";
			LineBuffer0(423) <= "00000000";
			LineBuffer0(424) <= "00000000";
			LineBuffer0(425) <= "00000000";
			LineBuffer0(426) <= "00000000";
			LineBuffer0(427) <= "00000000";
			LineBuffer0(428) <= "00000000";
			LineBuffer0(429) <= "00000000";	
			LineBuffer0(430) <= "00000000";
			LineBuffer0(431) <= "00000000";
			LineBuffer0(432) <= "00000000";
			LineBuffer0(433) <= "00000000";
			LineBuffer0(434) <= "00000000";
			LineBuffer0(435) <= "00000000";
			LineBuffer0(436) <= "00000000";
			LineBuffer0(437) <= "00000000";
			LineBuffer0(438) <= "00000000";
			LineBuffer0(439) <= "00000000";	
			LineBuffer0(440) <= "00000000";
			LineBuffer0(441) <= "00000000";
			LineBuffer0(442) <= "00000000";
			LineBuffer0(443) <= "00000000";
			LineBuffer0(444) <= "00000000";
			LineBuffer0(445) <= "00000000";
			LineBuffer0(446) <= "00000000";
			LineBuffer0(447) <= "00000000";
			LineBuffer0(448) <= "00000000";
			LineBuffer0(449) <= "00000000";	
			LineBuffer0(450) <= "00000000";
			LineBuffer0(451) <= "00000000";
			LineBuffer0(452) <= "00000000";
			LineBuffer0(453) <= "00000000";
			LineBuffer0(454) <= "00000000";
			LineBuffer0(455) <= "00000000";
			LineBuffer0(456) <= "00000000";
			LineBuffer0(457) <= "00000000";
			LineBuffer0(458) <= "00000000";
			LineBuffer0(459) <= "00000000";	
			LineBuffer0(460) <= "00000000";
			LineBuffer0(461) <= "00000000";
			LineBuffer0(462) <= "00000000";
			LineBuffer0(463) <= "00000000";
			LineBuffer0(464) <= "00000000";
			LineBuffer0(465) <= "00000000";
			LineBuffer0(466) <= "00000000";
			LineBuffer0(467) <= "00000000";
			LineBuffer0(468) <= "00000000";
			LineBuffer0(469) <= "00000000";	
			LineBuffer0(470) <= "00000000";
			LineBuffer0(471) <= "00000000";
			LineBuffer0(472) <= "00000000";
			LineBuffer0(473) <= "00000000";
			LineBuffer0(474) <= "00000000";
			LineBuffer0(475) <= "00000000";
			LineBuffer0(476) <= "00000000";
			LineBuffer0(477) <= "00000000";
			LineBuffer0(478) <= "00000000";
			LineBuffer0(479) <= "00000000";	
			LineBuffer0(480) <= "00000000";
			LineBuffer0(481) <= "00000000";
			LineBuffer0(482) <= "00000000";
			LineBuffer0(483) <= "00000000";
			LineBuffer0(484) <= "00000000";
			LineBuffer0(485) <= "00000000";
			LineBuffer0(486) <= "00000000";
			LineBuffer0(487) <= "00000000";
			LineBuffer0(488) <= "00000000";
			LineBuffer0(489) <= "00000000";	
			LineBuffer0(490) <= "00000000";
			LineBuffer0(491) <= "00000000";
			LineBuffer0(492) <= "00000000";
			LineBuffer0(493) <= "00000000";
			LineBuffer0(494) <= "00000000";
			LineBuffer0(495) <= "00000000";
			LineBuffer0(496) <= "00000000";
			LineBuffer0(497) <= "00000000";
			LineBuffer0(498) <= "00000000";
			LineBuffer0(499) <= "00000000";
			LineBuffer0(500) <= "00000000";
			LineBuffer0(501) <= "00000000";
			LineBuffer0(502) <= "00000000";
			LineBuffer0(503) <= "00000000";
			LineBuffer0(504) <= "00000000";
			LineBuffer0(505) <= "00000000";
			LineBuffer0(506) <= "00000000";
			LineBuffer0(507) <= "00000000";
			LineBuffer0(508) <= "00000000";
			LineBuffer0(509) <= "00000000";	
			LineBuffer0(510) <= "00000000";
			LineBuffer0(511) <= "00000000";
			LineBuffer0(512) <= "00000000";
			LineBuffer0(513) <= "00000000";
			LineBuffer0(514) <= "00000000";
			LineBuffer0(515) <= "00000000";
			LineBuffer0(516) <= "00000000";
			LineBuffer0(517) <= "00000000";
			LineBuffer0(518) <= "00000000";
			LineBuffer0(519) <= "00000000";	
			LineBuffer0(520) <= "00000000";
			LineBuffer0(521) <= "00000000";
			LineBuffer0(522) <= "00000000";
			LineBuffer0(523) <= "00000000";
			LineBuffer0(524) <= "00000000";
			LineBuffer0(525) <= "00000000";
			LineBuffer0(526) <= "00000000";
			LineBuffer0(527) <= "00000000";
			LineBuffer0(528) <= "00000000";
			LineBuffer0(529) <= "00000000";	
			LineBuffer0(530) <= "00000000";
			LineBuffer0(531) <= "00000000";
			LineBuffer0(532) <= "00000000";
			LineBuffer0(533) <= "00000000";
			LineBuffer0(534) <= "00000000";
			LineBuffer0(535) <= "00000000";
			LineBuffer0(536) <= "00000000";
			LineBuffer0(537) <= "00000000";
			LineBuffer0(538) <= "00000000";
			LineBuffer0(539) <= "00000000";	
			LineBuffer0(540) <= "00000000";
			LineBuffer0(541) <= "00000000";
			LineBuffer0(542) <= "00000000";
			LineBuffer0(543) <= "00000000";
			LineBuffer0(544) <= "00000000";
			LineBuffer0(545) <= "00000000";
			LineBuffer0(546) <= "00000000";
			LineBuffer0(547) <= "00000000";
			LineBuffer0(548) <= "00000000";
			LineBuffer0(549) <= "00000000";	
			LineBuffer0(550) <= "00000000";
			LineBuffer0(551) <= "00000000";
			LineBuffer0(552) <= "00000000";
			LineBuffer0(553) <= "00000000";
			LineBuffer0(554) <= "00000000";
			LineBuffer0(555) <= "00000000";
			LineBuffer0(556) <= "00000000";
			LineBuffer0(557) <= "00000000";
			LineBuffer0(558) <= "00000000";
			LineBuffer0(559) <= "00000000";	
			LineBuffer0(560) <= "00000000";
			LineBuffer0(561) <= "00000000";
			LineBuffer0(562) <= "00000000";
			LineBuffer0(563) <= "00000000";
			LineBuffer0(564) <= "00000000";
			LineBuffer0(565) <= "00000000";
			LineBuffer0(566) <= "00000000";
			LineBuffer0(567) <= "00000000";
			LineBuffer0(568) <= "00000000";
			LineBuffer0(569) <= "00000000";	
			LineBuffer0(570) <= "00000000";
			LineBuffer0(571) <= "00000000";
			LineBuffer0(572) <= "00000000";
			LineBuffer0(573) <= "00000000";
			LineBuffer0(574) <= "00000000";
			LineBuffer0(575) <= "00000000";
			LineBuffer0(576) <= "00000000";
			LineBuffer0(577) <= "00000000";
			LineBuffer0(578) <= "00000000";
			LineBuffer0(579) <= "00000000";	
			LineBuffer0(580) <= "00000000";
			LineBuffer0(581) <= "00000000";
			LineBuffer0(582) <= "00000000";
			LineBuffer0(583) <= "00000000";
			LineBuffer0(584) <= "00000000";
			LineBuffer0(585) <= "00000000";
			LineBuffer0(586) <= "00000000";
			LineBuffer0(587) <= "00000000";
			LineBuffer0(588) <= "00000000";
			LineBuffer0(589) <= "00000000";	
			LineBuffer0(590) <= "00000000";
			LineBuffer0(591) <= "00000000";
			LineBuffer0(592) <= "00000000";
			LineBuffer0(593) <= "00000000";
			LineBuffer0(594) <= "00000000";
			LineBuffer0(595) <= "00000000";
			LineBuffer0(596) <= "00000000";
			LineBuffer0(597) <= "00000000";
			LineBuffer0(598) <= "00000000";
			LineBuffer0(599) <= "00000000";
			LineBuffer0(600) <= "00000000";
			LineBuffer0(601) <= "00000000";
			LineBuffer0(602) <= "00000000";
			LineBuffer0(603) <= "00000000";
			LineBuffer0(604) <= "00000000";
			LineBuffer0(605) <= "00000000";
			LineBuffer0(606) <= "00000000";
			LineBuffer0(607) <= "00000000";
			LineBuffer0(608) <= "00000000";
			LineBuffer0(609) <= "00000000";	
			LineBuffer0(610) <= "00000000";
			LineBuffer0(611) <= "00000000";
			LineBuffer0(612) <= "00000000";
			LineBuffer0(613) <= "00000000";
			LineBuffer0(614) <= "00000000";
			LineBuffer0(615) <= "00000000";
			LineBuffer0(616) <= "00000000";
			LineBuffer0(617) <= "00000000";
			LineBuffer0(618) <= "00000000";
			LineBuffer0(619) <= "00000000";	
			LineBuffer0(620) <= "00000000";
			LineBuffer0(621) <= "00000000";
			LineBuffer0(622) <= "00000000";
			LineBuffer0(623) <= "00000000";
			LineBuffer0(624) <= "00000000";
			LineBuffer0(625) <= "00000000";
			LineBuffer0(626) <= "00000000";
			LineBuffer0(627) <= "00000000";
			LineBuffer0(628) <= "00000000";
			LineBuffer0(629) <= "00000000";	
			LineBuffer0(630) <= "00000000";
			LineBuffer0(631) <= "00000000";
			LineBuffer0(632) <= "00000000";
			LineBuffer0(633) <= "00000000";
			LineBuffer0(634) <= "00000000";
			LineBuffer0(635) <= "00000000";
			LineBuffer0(636) <= "00000000";
			LineBuffer0(637) <= "00000000";
			LineBuffer0(638) <= "00000000";
			LineBuffer0(639) <= "00000000";
			LineBuffer0(640) <= "00000000";
            LineBuffer0(641) <= "00000000";
            LineBuffer0(642) <= "00000000";
            LineBuffer0(643) <= "00000000";
            LineBuffer0(644) <= "00000000";
            LineBuffer0(645) <= "00000000";
            LineBuffer0(646) <= "00000000";
            LineBuffer0(647) <= "00000000";
            LineBuffer0(648) <= "00000000";
            LineBuffer0(649) <= "00000000";    
            LineBuffer0(650) <= "00000000";
            LineBuffer0(651) <= "00000000";
            LineBuffer0(652) <= "00000000";
            LineBuffer0(653) <= "00000000";
            LineBuffer0(654) <= "00000000";
            LineBuffer0(655) <= "00000000";
            LineBuffer0(656) <= "00000000";
            LineBuffer0(657) <= "00000000";
            LineBuffer0(658) <= "00000000";
            LineBuffer0(659) <= "00000000";    
            LineBuffer0(660) <= "00000000";
            LineBuffer0(661) <= "00000000";
            LineBuffer0(662) <= "00000000";
            LineBuffer0(663) <= "00000000";
            LineBuffer0(664) <= "00000000";
            LineBuffer0(665) <= "00000000";
            LineBuffer0(666) <= "00000000";
            LineBuffer0(667) <= "00000000";
            LineBuffer0(668) <= "00000000";
            LineBuffer0(669) <= "00000000";    
            LineBuffer0(670) <= "00000000";
            LineBuffer0(671) <= "00000000";
            LineBuffer0(672) <= "00000000";
            LineBuffer0(673) <= "00000000";
            LineBuffer0(674) <= "00000000";
            LineBuffer0(675) <= "00000000";
            LineBuffer0(676) <= "00000000";
            LineBuffer0(677) <= "00000000";
            LineBuffer0(678) <= "00000000";
            LineBuffer0(679) <= "00000000";    
            LineBuffer0(680) <= "00000000";
            LineBuffer0(681) <= "00000000";
            LineBuffer0(682) <= "00000000";
            LineBuffer0(683) <= "00000000";
            LineBuffer0(684) <= "00000000";
            LineBuffer0(685) <= "00000000";
            LineBuffer0(686) <= "00000000";
            LineBuffer0(687) <= "00000000";
            LineBuffer0(688) <= "00000000";
            LineBuffer0(689) <= "00000000";    
            LineBuffer0(690) <= "00000000";
            LineBuffer0(691) <= "00000000";
            LineBuffer0(692) <= "00000000";
            LineBuffer0(693) <= "00000000";
            LineBuffer0(694) <= "00000000";
            LineBuffer0(695) <= "00000000";
            LineBuffer0(696) <= "00000000";
            LineBuffer0(697) <= "00000000";
            LineBuffer0(698) <= "00000000";
            LineBuffer0(699) <= "00000000";    
            LineBuffer0(700) <= "00000000";
            LineBuffer0(701) <= "00000000";
            LineBuffer0(702) <= "00000000";
            LineBuffer0(703) <= "00000000";
            LineBuffer0(704) <= "00000000";
            LineBuffer0(705) <= "00000000";
            LineBuffer0(706) <= "00000000";
            LineBuffer0(707) <= "00000000";
            LineBuffer0(708) <= "00000000";
            LineBuffer0(709) <= "00000000";    
            LineBuffer0(710) <= "00000000";
            LineBuffer0(711) <= "00000000";
            LineBuffer0(712) <= "00000000";
            LineBuffer0(713) <= "00000000";
            LineBuffer0(714) <= "00000000";
            LineBuffer0(715) <= "00000000";
            LineBuffer0(716) <= "00000000";
            LineBuffer0(717) <= "00000000";
            LineBuffer0(718) <= "00000000";
            LineBuffer0(719) <= "00000000";    
            LineBuffer0(720) <= "00000000";
            LineBuffer0(721) <= "00000000";
            LineBuffer0(722) <= "00000000";
            LineBuffer0(723) <= "00000000";
            LineBuffer0(724) <= "00000000";
            LineBuffer0(725) <= "00000000";
            LineBuffer0(726) <= "00000000";
            LineBuffer0(727) <= "00000000";
            LineBuffer0(728) <= "00000000";
            LineBuffer0(729) <= "00000000";    
            LineBuffer0(730) <= "00000000";
            LineBuffer0(731) <= "00000000";
            LineBuffer0(732) <= "00000000";
            LineBuffer0(733) <= "00000000";
            LineBuffer0(734) <= "00000000";
            LineBuffer0(735) <= "00000000";
            LineBuffer0(736) <= "00000000";
            LineBuffer0(737) <= "00000000";
            LineBuffer0(738) <= "00000000";
            LineBuffer0(739) <= "00000000";    
            LineBuffer0(740) <= "00000000";
            LineBuffer0(741) <= "00000000";
            LineBuffer0(742) <= "00000000";
            LineBuffer0(743) <= "00000000";
            LineBuffer0(744) <= "00000000";
            LineBuffer0(745) <= "00000000";
            LineBuffer0(746) <= "00000000";
            LineBuffer0(747) <= "00000000";
            LineBuffer0(748) <= "00000000";
            LineBuffer0(749) <= "00000000";    
            LineBuffer0(750) <= "00000000";
            LineBuffer0(751) <= "00000000";
            LineBuffer0(752) <= "00000000";
            LineBuffer0(753) <= "00000000";
            LineBuffer0(754) <= "00000000";
            LineBuffer0(755) <= "00000000";
            LineBuffer0(756) <= "00000000";
            LineBuffer0(757) <= "00000000";
            LineBuffer0(758) <= "00000000";
            LineBuffer0(759) <= "00000000";    
            LineBuffer0(760) <= "00000000";
            LineBuffer0(761) <= "00000000";
            LineBuffer0(762) <= "00000000";
            LineBuffer0(763) <= "00000000";
            LineBuffer0(764) <= "00000000";
            LineBuffer0(765) <= "00000000";
            LineBuffer0(766) <= "00000000";
            LineBuffer0(767) <= "00000000";
            LineBuffer0(768) <= "00000000";
            LineBuffer0(769) <= "00000000";    
            LineBuffer0(770) <= "00000000";
            LineBuffer0(771) <= "00000000";
            LineBuffer0(772) <= "00000000";
            LineBuffer0(773) <= "00000000";
            LineBuffer0(774) <= "00000000";
            LineBuffer0(775) <= "00000000";
            LineBuffer0(776) <= "00000000";
            LineBuffer0(777) <= "00000000";
            LineBuffer0(778) <= "00000000";
            LineBuffer0(779) <= "00000000";    
            LineBuffer0(780) <= "00000000";
            LineBuffer0(781) <= "00000000";
            LineBuffer0(782) <= "00000000";
            LineBuffer0(783) <= "00000000";
            LineBuffer0(784) <= "00000000";
            LineBuffer0(785) <= "00000000";
            LineBuffer0(786) <= "00000000";
            LineBuffer0(787) <= "00000000";
            LineBuffer0(788) <= "00000000";
            LineBuffer0(789) <= "00000000";    
            LineBuffer0(790) <= "00000000";
            LineBuffer0(791) <= "00000000";
            LineBuffer0(792) <= "00000000";
            LineBuffer0(793) <= "00000000";
            LineBuffer0(794) <= "00000000";
            LineBuffer0(795) <= "00000000";
            LineBuffer0(796) <= "00000000";
            LineBuffer0(797) <= "00000000";
            LineBuffer0(798) <= "00000000";
            LineBuffer0(799) <= "00000000";    
            LineBuffer0(800) <= "00000000";
            LineBuffer0(801) <= "00000000";
            LineBuffer0(802) <= "00000000";
            LineBuffer0(803) <= "00000000";
            LineBuffer0(804) <= "00000000";
            LineBuffer0(805) <= "00000000";
            LineBuffer0(806) <= "00000000";
            LineBuffer0(807) <= "00000000";
            LineBuffer0(808) <= "00000000";
            LineBuffer0(809) <= "00000000";    
            LineBuffer0(810) <= "00000000";
            LineBuffer0(811) <= "00000000";
            LineBuffer0(812) <= "00000000";
            LineBuffer0(813) <= "00000000";
            LineBuffer0(814) <= "00000000";
            LineBuffer0(815) <= "00000000";
            LineBuffer0(816) <= "00000000";
            LineBuffer0(817) <= "00000000";
            LineBuffer0(818) <= "00000000";
            LineBuffer0(819) <= "00000000";    
            LineBuffer0(820) <= "00000000";
            LineBuffer0(821) <= "00000000";
            LineBuffer0(822) <= "00000000";
            LineBuffer0(823) <= "00000000";
            LineBuffer0(824) <= "00000000";
            LineBuffer0(825) <= "00000000";
            LineBuffer0(826) <= "00000000";
            LineBuffer0(827) <= "00000000";
            LineBuffer0(828) <= "00000000";
            LineBuffer0(829) <= "00000000";    
            LineBuffer0(830) <= "00000000";
            LineBuffer0(831) <= "00000000";
            LineBuffer0(832) <= "00000000";
            LineBuffer0(833) <= "00000000";
            LineBuffer0(834) <= "00000000";
            LineBuffer0(835) <= "00000000";
            LineBuffer0(836) <= "00000000";
            LineBuffer0(837) <= "00000000";
            LineBuffer0(838) <= "00000000";
            LineBuffer0(839) <= "00000000";
            LineBuffer0(840) <= "00000000";
            LineBuffer0(841) <= "00000000";
            LineBuffer0(842) <= "00000000";
            LineBuffer0(843) <= "00000000";
            LineBuffer0(844) <= "00000000";
            LineBuffer0(845) <= "00000000";
            LineBuffer0(846) <= "00000000";
            LineBuffer0(847) <= "00000000";
            LineBuffer0(848) <= "00000000";
            LineBuffer0(849) <= "00000000";    
            LineBuffer0(850) <= "00000000";
            LineBuffer0(851) <= "00000000";
            LineBuffer0(852) <= "00000000";
            LineBuffer0(853) <= "00000000";
            LineBuffer0(854) <= "00000000";
            LineBuffer0(855) <= "00000000";
            LineBuffer0(856) <= "00000000";
            LineBuffer0(857) <= "00000000";
            LineBuffer0(858) <= "00000000";
            LineBuffer0(859) <= "00000000";    
            LineBuffer0(860) <= "00000000";
            LineBuffer0(861) <= "00000000";
            LineBuffer0(862) <= "00000000";
            LineBuffer0(863) <= "00000000";
            LineBuffer0(864) <= "00000000";
            LineBuffer0(865) <= "00000000";
            LineBuffer0(866) <= "00000000";
            LineBuffer0(867) <= "00000000";
            LineBuffer0(868) <= "00000000";
            LineBuffer0(869) <= "00000000";    
            LineBuffer0(870) <= "00000000";
            LineBuffer0(871) <= "00000000";
            LineBuffer0(872) <= "00000000";
            LineBuffer0(873) <= "00000000";
            LineBuffer0(874) <= "00000000";
            LineBuffer0(875) <= "00000000";
            LineBuffer0(876) <= "00000000";
            LineBuffer0(877) <= "00000000";
            LineBuffer0(878) <= "00000000";
            LineBuffer0(879) <= "00000000";    
            LineBuffer0(880) <= "00000000";
            LineBuffer0(881) <= "00000000";
            LineBuffer0(882) <= "00000000";
            LineBuffer0(883) <= "00000000";
            LineBuffer0(884) <= "00000000";
            LineBuffer0(885) <= "00000000";
            LineBuffer0(886) <= "00000000";
            LineBuffer0(887) <= "00000000";
            LineBuffer0(888) <= "00000000";
            LineBuffer0(889) <= "00000000";    
            LineBuffer0(890) <= "00000000";
            LineBuffer0(891) <= "00000000";
            LineBuffer0(892) <= "00000000";
            LineBuffer0(893) <= "00000000";
            LineBuffer0(894) <= "00000000";
            LineBuffer0(895) <= "00000000";
            LineBuffer0(896) <= "00000000";
            LineBuffer0(897) <= "00000000";
            LineBuffer0(898) <= "00000000";
            LineBuffer0(899) <= "00000000";    
            LineBuffer0(900) <= "00000000";
            LineBuffer0(901) <= "00000000";
            LineBuffer0(902) <= "00000000";
            LineBuffer0(903) <= "00000000";
            LineBuffer0(904) <= "00000000";
            LineBuffer0(905) <= "00000000";
            LineBuffer0(906) <= "00000000";
            LineBuffer0(907) <= "00000000";
            LineBuffer0(908) <= "00000000";
            LineBuffer0(909) <= "00000000";    
            LineBuffer0(910) <= "00000000";
            LineBuffer0(911) <= "00000000";
            LineBuffer0(912) <= "00000000";
            LineBuffer0(913) <= "00000000";
            LineBuffer0(914) <= "00000000";
            LineBuffer0(915) <= "00000000";
            LineBuffer0(916) <= "00000000";
            LineBuffer0(917) <= "00000000";
            LineBuffer0(918) <= "00000000";
            LineBuffer0(919) <= "00000000";    
            LineBuffer0(920) <= "00000000";
            LineBuffer0(921) <= "00000000";
            LineBuffer0(922) <= "00000000";
            LineBuffer0(923) <= "00000000";
            LineBuffer0(924) <= "00000000";
            LineBuffer0(925) <= "00000000";
            LineBuffer0(926) <= "00000000";
            LineBuffer0(927) <= "00000000";
            LineBuffer0(928) <= "00000000";
            LineBuffer0(929) <= "00000000";    
            LineBuffer0(930) <= "00000000";
            LineBuffer0(931) <= "00000000";
            LineBuffer0(932) <= "00000000";
            LineBuffer0(933) <= "00000000";
            LineBuffer0(934) <= "00000000";
            LineBuffer0(935) <= "00000000";
            LineBuffer0(936) <= "00000000";
            LineBuffer0(937) <= "00000000";
            LineBuffer0(938) <= "00000000";
            LineBuffer0(939) <= "00000000";
            LineBuffer0(940) <= "00000000";
            LineBuffer0(941) <= "00000000";
            LineBuffer0(942) <= "00000000";
            LineBuffer0(943) <= "00000000";
            LineBuffer0(944) <= "00000000";
            LineBuffer0(945) <= "00000000";
            LineBuffer0(946) <= "00000000";
            LineBuffer0(947) <= "00000000";
            LineBuffer0(948) <= "00000000";
            LineBuffer0(949) <= "00000000";    
            LineBuffer0(950) <= "00000000";
            LineBuffer0(951) <= "00000000";
            LineBuffer0(952) <= "00000000";
            LineBuffer0(953) <= "00000000";
            LineBuffer0(954) <= "00000000";
            LineBuffer0(955) <= "00000000";
            LineBuffer0(956) <= "00000000";
            LineBuffer0(957) <= "00000000";
            LineBuffer0(958) <= "00000000";
            LineBuffer0(959) <= "00000000";    
            LineBuffer0(960) <= "00000000";
            LineBuffer0(961) <= "00000000";
            LineBuffer0(962) <= "00000000";
            LineBuffer0(963) <= "00000000";
            LineBuffer0(964) <= "00000000";
            LineBuffer0(965) <= "00000000";
            LineBuffer0(966) <= "00000000";
            LineBuffer0(967) <= "00000000";
            LineBuffer0(968) <= "00000000";
            LineBuffer0(969) <= "00000000";    
            LineBuffer0(970) <= "00000000";
            LineBuffer0(971) <= "00000000";
            LineBuffer0(972) <= "00000000";
            LineBuffer0(973) <= "00000000";
            LineBuffer0(974) <= "00000000";
            LineBuffer0(975) <= "00000000";
            LineBuffer0(976) <= "00000000";
            LineBuffer0(977) <= "00000000";
            LineBuffer0(978) <= "00000000";
            LineBuffer0(979) <= "00000000";    
            LineBuffer0(980) <= "00000000";
            LineBuffer0(981) <= "00000000";
            LineBuffer0(982) <= "00000000";
            LineBuffer0(983) <= "00000000";
            LineBuffer0(984) <= "00000000";
            LineBuffer0(985) <= "00000000";
            LineBuffer0(986) <= "00000000";
            LineBuffer0(987) <= "00000000";
            LineBuffer0(988) <= "00000000";
            LineBuffer0(989) <= "00000000";    
            LineBuffer0(990) <= "00000000";
            LineBuffer0(991) <= "00000000";
            LineBuffer0(992) <= "00000000";
            LineBuffer0(993) <= "00000000";
            LineBuffer0(994) <= "00000000";
            LineBuffer0(995) <= "00000000";
            LineBuffer0(996) <= "00000000";
            LineBuffer0(997) <= "00000000";
            LineBuffer0(998) <= "00000000";
            LineBuffer0(999) <= "00000000";    
            LineBuffer0(1000) <= "00000000";
            LineBuffer0(1001) <= "00000000";
            LineBuffer0(1002) <= "00000000";
            LineBuffer0(1003) <= "00000000";
            LineBuffer0(1004) <= "00000000";
            LineBuffer0(1005) <= "00000000";
            LineBuffer0(1006) <= "00000000";
            LineBuffer0(1007) <= "00000000";
            LineBuffer0(1008) <= "00000000";
            LineBuffer0(1009) <= "00000000";    
            LineBuffer0(1010) <= "00000000";
            LineBuffer0(1011) <= "00000000";
            LineBuffer0(1012) <= "00000000";
            LineBuffer0(1013) <= "00000000";
            LineBuffer0(1014) <= "00000000";
            LineBuffer0(1015) <= "00000000";
            LineBuffer0(1016) <= "00000000";
            LineBuffer0(1017) <= "00000000";
            LineBuffer0(1018) <= "00000000";
            LineBuffer0(1019) <= "00000000";    
            LineBuffer0(1020) <= "00000000";
            LineBuffer0(1021) <= "00000000";
            LineBuffer0(1022) <= "00000000";
            LineBuffer0(1023) <= "00000000";
            LineBuffer0(1024) <= "00000000";
            LineBuffer0(1025) <= "00000000";
            LineBuffer0(1026) <= "00000000";
            LineBuffer0(1027) <= "00000000";
            LineBuffer0(1028) <= "00000000";
            LineBuffer0(1029) <= "00000000";    
            LineBuffer0(1030) <= "00000000";
            LineBuffer0(1031) <= "00000000";
            LineBuffer0(1032) <= "00000000";
            LineBuffer0(1033) <= "00000000";
            LineBuffer0(1034) <= "00000000";
            LineBuffer0(1035) <= "00000000";
            LineBuffer0(1036) <= "00000000";
            LineBuffer0(1037) <= "00000000";
            LineBuffer0(1038) <= "00000000";
            LineBuffer0(1039) <= "00000000";
            LineBuffer0(1040) <= "00000000";
            LineBuffer0(1041) <= "00000000";
            LineBuffer0(1042) <= "00000000";
            LineBuffer0(1043) <= "00000000";
            LineBuffer0(1044) <= "00000000";
            LineBuffer0(1045) <= "00000000";
            LineBuffer0(1046) <= "00000000";
            LineBuffer0(1047) <= "00000000";
            LineBuffer0(1048) <= "00000000";
            LineBuffer0(1049) <= "00000000";    
            LineBuffer0(1050) <= "00000000";
            LineBuffer0(1051) <= "00000000";
            LineBuffer0(1052) <= "00000000";
            LineBuffer0(1053) <= "00000000";
            LineBuffer0(1054) <= "00000000";
            LineBuffer0(1055) <= "00000000";
            LineBuffer0(1056) <= "00000000";
            LineBuffer0(1057) <= "00000000";
            LineBuffer0(1058) <= "00000000";
            LineBuffer0(1059) <= "00000000";    
            LineBuffer0(1060) <= "00000000";
            LineBuffer0(1061) <= "00000000";
            LineBuffer0(1062) <= "00000000";
            LineBuffer0(1063) <= "00000000";
            LineBuffer0(1064) <= "00000000";
            LineBuffer0(1065) <= "00000000";
            LineBuffer0(1066) <= "00000000";
            LineBuffer0(1067) <= "00000000";
            LineBuffer0(1068) <= "00000000";
            LineBuffer0(1069) <= "00000000";    
            LineBuffer0(1070) <= "00000000";
            LineBuffer0(1071) <= "00000000";
            LineBuffer0(1072) <= "00000000";
            LineBuffer0(1073) <= "00000000";
            LineBuffer0(1074) <= "00000000";
            LineBuffer0(1075) <= "00000000";
            LineBuffer0(1076) <= "00000000";
            LineBuffer0(1077) <= "00000000";
            LineBuffer0(1078) <= "00000000";
            LineBuffer0(1079) <= "00000000";    
            LineBuffer0(1080) <= "00000000";
            LineBuffer0(1081) <= "00000000";
            LineBuffer0(1082) <= "00000000";
            LineBuffer0(1083) <= "00000000";
            LineBuffer0(1084) <= "00000000";
            LineBuffer0(1085) <= "00000000";
            LineBuffer0(1086) <= "00000000";
            LineBuffer0(1087) <= "00000000";
            LineBuffer0(1088) <= "00000000";
            LineBuffer0(1089) <= "00000000";    
            LineBuffer0(1090) <= "00000000";
            LineBuffer0(1091) <= "00000000";
            LineBuffer0(1092) <= "00000000";
            LineBuffer0(1093) <= "00000000";
            LineBuffer0(1094) <= "00000000";
            LineBuffer0(1095) <= "00000000";
            LineBuffer0(1096) <= "00000000";
            LineBuffer0(1097) <= "00000000";
            LineBuffer0(1098) <= "00000000";
            LineBuffer0(1099) <= "00000000";    
            LineBuffer0(1100) <= "00000000";
            LineBuffer0(1101) <= "00000000";
            LineBuffer0(1102) <= "00000000";
            LineBuffer0(1103) <= "00000000";
            LineBuffer0(1104) <= "00000000";
            LineBuffer0(1105) <= "00000000";
            LineBuffer0(1106) <= "00000000";
            LineBuffer0(1107) <= "00000000";
            LineBuffer0(1108) <= "00000000";
            LineBuffer0(1109) <= "00000000";    
            LineBuffer0(1110) <= "00000000";
            LineBuffer0(1111) <= "00000000";
            LineBuffer0(1112) <= "00000000";
            LineBuffer0(1113) <= "00000000";
            LineBuffer0(1114) <= "00000000";
            LineBuffer0(1115) <= "00000000";
            LineBuffer0(1116) <= "00000000";
            LineBuffer0(1117) <= "00000000";
            LineBuffer0(1118) <= "00000000";
            LineBuffer0(1119) <= "00000000";    
            LineBuffer0(1120) <= "00000000";
            LineBuffer0(1121) <= "00000000";
            LineBuffer0(1122) <= "00000000";
            LineBuffer0(1123) <= "00000000";
            LineBuffer0(1124) <= "00000000";
            LineBuffer0(1125) <= "00000000";
            LineBuffer0(1126) <= "00000000";
            LineBuffer0(1127) <= "00000000";
            LineBuffer0(1128) <= "00000000";
            LineBuffer0(1129) <= "00000000";    
            LineBuffer0(1130) <= "00000000";
            LineBuffer0(1131) <= "00000000";
            LineBuffer0(1132) <= "00000000";
            LineBuffer0(1133) <= "00000000";
            LineBuffer0(1134) <= "00000000";
            LineBuffer0(1135) <= "00000000";
            LineBuffer0(1136) <= "00000000";
            LineBuffer0(1137) <= "00000000";
            LineBuffer0(1138) <= "00000000";
            LineBuffer0(1139) <= "00000000";
            LineBuffer0(1140) <= "00000000";
            LineBuffer0(1141) <= "00000000";
            LineBuffer0(1142) <= "00000000";
            LineBuffer0(1143) <= "00000000";
            LineBuffer0(1144) <= "00000000";
            LineBuffer0(1145) <= "00000000";
            LineBuffer0(1146) <= "00000000";
            LineBuffer0(1147) <= "00000000";
            LineBuffer0(1148) <= "00000000";
            LineBuffer0(1149) <= "00000000";    
            LineBuffer0(1150) <= "00000000";
            LineBuffer0(1151) <= "00000000";
            LineBuffer0(1152) <= "00000000";
            LineBuffer0(1153) <= "00000000";
            LineBuffer0(1154) <= "00000000";
            LineBuffer0(1155) <= "00000000";
            LineBuffer0(1156) <= "00000000";
            LineBuffer0(1157) <= "00000000";
            LineBuffer0(1158) <= "00000000";
            LineBuffer0(1159) <= "00000000";    
            LineBuffer0(1160) <= "00000000";
            LineBuffer0(1161) <= "00000000";
            LineBuffer0(1162) <= "00000000";
            LineBuffer0(1163) <= "00000000";
            LineBuffer0(1164) <= "00000000";
            LineBuffer0(1165) <= "00000000";
            LineBuffer0(1166) <= "00000000";
            LineBuffer0(1167) <= "00000000";
            LineBuffer0(1168) <= "00000000";
            LineBuffer0(1169) <= "00000000";    
            LineBuffer0(1170) <= "00000000";
            LineBuffer0(1171) <= "00000000";
            LineBuffer0(1172) <= "00000000";
            LineBuffer0(1173) <= "00000000";
            LineBuffer0(1174) <= "00000000";
            LineBuffer0(1175) <= "00000000";
            LineBuffer0(1176) <= "00000000";
            LineBuffer0(1177) <= "00000000";
            LineBuffer0(1178) <= "00000000";
            LineBuffer0(1179) <= "00000000";    
            LineBuffer0(1180) <= "00000000";
            LineBuffer0(1181) <= "00000000";
            LineBuffer0(1182) <= "00000000";
            LineBuffer0(1183) <= "00000000";
            LineBuffer0(1184) <= "00000000";
            LineBuffer0(1185) <= "00000000";
            LineBuffer0(1186) <= "00000000";
            LineBuffer0(1187) <= "00000000";
            LineBuffer0(1188) <= "00000000";
            LineBuffer0(1189) <= "00000000";    
            LineBuffer0(1190) <= "00000000";
            LineBuffer0(1191) <= "00000000";
            LineBuffer0(1192) <= "00000000";
            LineBuffer0(1193) <= "00000000";
            LineBuffer0(1194) <= "00000000";
            LineBuffer0(1195) <= "00000000";
            LineBuffer0(1196) <= "00000000";
            LineBuffer0(1197) <= "00000000";
            LineBuffer0(1198) <= "00000000";
            LineBuffer0(1199) <= "00000000";    
            LineBuffer0(1200) <= "00000000";
            LineBuffer0(1201) <= "00000000";
            LineBuffer0(1202) <= "00000000";
            LineBuffer0(1203) <= "00000000";
            LineBuffer0(1204) <= "00000000";
            LineBuffer0(1205) <= "00000000";
            LineBuffer0(1206) <= "00000000";
            LineBuffer0(1207) <= "00000000";
            LineBuffer0(1208) <= "00000000";
            LineBuffer0(1209) <= "00000000";    
            LineBuffer0(1210) <= "00000000";
            LineBuffer0(1211) <= "00000000";
            LineBuffer0(1212) <= "00000000";
            LineBuffer0(1213) <= "00000000";
            LineBuffer0(1214) <= "00000000";
            LineBuffer0(1215) <= "00000000";
            LineBuffer0(1216) <= "00000000";
            LineBuffer0(1217) <= "00000000";
            LineBuffer0(1218) <= "00000000";
            LineBuffer0(1219) <= "00000000";    
            LineBuffer0(1220) <= "00000000";
            LineBuffer0(1221) <= "00000000";
            LineBuffer0(1222) <= "00000000";
            LineBuffer0(1223) <= "00000000";
            LineBuffer0(1224) <= "00000000";
            LineBuffer0(1225) <= "00000000";
            LineBuffer0(1226) <= "00000000";
            LineBuffer0(1227) <= "00000000";
            LineBuffer0(1228) <= "00000000";
            LineBuffer0(1229) <= "00000000";    
            LineBuffer0(1230) <= "00000000";
            LineBuffer0(1231) <= "00000000";
            LineBuffer0(1232) <= "00000000";
            LineBuffer0(1233) <= "00000000";
            LineBuffer0(1234) <= "00000000";
            LineBuffer0(1235) <= "00000000";
            LineBuffer0(1236) <= "00000000";
            LineBuffer0(1237) <= "00000000";
            LineBuffer0(1238) <= "00000000";
            LineBuffer0(1239) <= "00000000";
            LineBuffer0(1240) <= "00000000";
            LineBuffer0(1241) <= "00000000";
            LineBuffer0(1242) <= "00000000";
            LineBuffer0(1243) <= "00000000";
            LineBuffer0(1244) <= "00000000";
            LineBuffer0(1245) <= "00000000";
            LineBuffer0(1246) <= "00000000";
            LineBuffer0(1247) <= "00000000";
            LineBuffer0(1248) <= "00000000";
            LineBuffer0(1249) <= "00000000";    
            LineBuffer0(1250) <= "00000000";
            LineBuffer0(1251) <= "00000000";
            LineBuffer0(1252) <= "00000000";
            LineBuffer0(1253) <= "00000000";
            LineBuffer0(1254) <= "00000000";
            LineBuffer0(1255) <= "00000000";
            LineBuffer0(1256) <= "00000000";
            LineBuffer0(1257) <= "00000000";
            LineBuffer0(1258) <= "00000000";
            LineBuffer0(1259) <= "00000000";    
            LineBuffer0(1260) <= "00000000";
            LineBuffer0(1261) <= "00000000";
            LineBuffer0(1262) <= "00000000";
            LineBuffer0(1263) <= "00000000";
            LineBuffer0(1264) <= "00000000";
            LineBuffer0(1265) <= "00000000";
            LineBuffer0(1266) <= "00000000";
            LineBuffer0(1267) <= "00000000";
            LineBuffer0(1268) <= "00000000";
            LineBuffer0(1269) <= "00000000";    
            LineBuffer0(1270) <= "00000000";
            LineBuffer0(1271) <= "00000000";
            LineBuffer0(1272) <= "00000000";
            LineBuffer0(1273) <= "00000000";
            LineBuffer0(1274) <= "00000000";
            LineBuffer0(1275) <= "00000000";
            LineBuffer0(1276) <= "00000000";
            LineBuffer0(1277) <= "00000000";
            LineBuffer0(1278) <= "00000000";
            LineBuffer0(1279) <= "00000000";
            
--			LineBuffer0(1280) <= "00000000";
--            LineBuffer0(1281) <= "00000000";
--            LineBuffer0(1282) <= "00000000";
--            LineBuffer0(1283) <= "00000000";
--            LineBuffer0(1284) <= "00000000";
--            LineBuffer0(1285) <= "00000000";
--            LineBuffer0(1286) <= "00000000";
--            LineBuffer0(1287) <= "00000000";
--            LineBuffer0(1288) <= "00000000";
--            LineBuffer0(1289) <= "00000000";    
--            LineBuffer0(1290) <= "00000000";
--            LineBuffer0(1291) <= "00000000";
--            LineBuffer0(1292) <= "00000000";
--            LineBuffer0(1293) <= "00000000";
--            LineBuffer0(1294) <= "00000000";
--            LineBuffer0(1295) <= "00000000";
--            LineBuffer0(1296) <= "00000000";
--            LineBuffer0(1297) <= "00000000";
--            LineBuffer0(1298) <= "00000000";
--            LineBuffer0(1299) <= "00000000";    
--            LineBuffer0(1300) <= "00000000";
--            LineBuffer0(1301) <= "00000000";
--            LineBuffer0(1302) <= "00000000";
--            LineBuffer0(1303) <= "00000000";
--            LineBuffer0(1304) <= "00000000";
--            LineBuffer0(1305) <= "00000000";
--            LineBuffer0(1306) <= "00000000";
--            LineBuffer0(1307) <= "00000000";
--            LineBuffer0(1308) <= "00000000";
--            LineBuffer0(1309) <= "00000000";    
--            LineBuffer0(1310) <= "00000000";
--            LineBuffer0(1311) <= "00000000";
--            LineBuffer0(1312) <= "00000000";
--            LineBuffer0(1313) <= "00000000";
--            LineBuffer0(1314) <= "00000000";
--            LineBuffer0(1315) <= "00000000";
--            LineBuffer0(1316) <= "00000000";
--            LineBuffer0(1317) <= "00000000";
--            LineBuffer0(1318) <= "00000000";
--            LineBuffer0(1319) <= "00000000";    
--            LineBuffer0(1320) <= "00000000";
--            LineBuffer0(1321) <= "00000000";
--            LineBuffer0(1322) <= "00000000";
--            LineBuffer0(1323) <= "00000000";
--            LineBuffer0(1324) <= "00000000";
--            LineBuffer0(1325) <= "00000000";
--            LineBuffer0(1326) <= "00000000";
--            LineBuffer0(1327) <= "00000000";
--            LineBuffer0(1328) <= "00000000";
--            LineBuffer0(1329) <= "00000000";    
--            LineBuffer0(1330) <= "00000000";
--            LineBuffer0(1331) <= "00000000";
--            LineBuffer0(1332) <= "00000000";
--            LineBuffer0(1333) <= "00000000";
--            LineBuffer0(1334) <= "00000000";
--            LineBuffer0(1335) <= "00000000";
--            LineBuffer0(1336) <= "00000000";
--            LineBuffer0(1337) <= "00000000";
--            LineBuffer0(1338) <= "00000000";
--            LineBuffer0(1339) <= "00000000";    
--            LineBuffer0(1340) <= "00000000";
--            LineBuffer0(1341) <= "00000000";
--            LineBuffer0(1342) <= "00000000";
--            LineBuffer0(1343) <= "00000000";
--            LineBuffer0(1344) <= "00000000";
--            LineBuffer0(1345) <= "00000000";
--            LineBuffer0(1346) <= "00000000";
--            LineBuffer0(1347) <= "00000000";
--            LineBuffer0(1348) <= "00000000";
--            LineBuffer0(1349) <= "00000000";    
--            LineBuffer0(1350) <= "00000000";
--            LineBuffer0(1351) <= "00000000";
--            LineBuffer0(1352) <= "00000000";
--            LineBuffer0(1353) <= "00000000";
--            LineBuffer0(1354) <= "00000000";
--            LineBuffer0(1355) <= "00000000";
--            LineBuffer0(1356) <= "00000000";
--            LineBuffer0(1357) <= "00000000";
--            LineBuffer0(1358) <= "00000000";
--            LineBuffer0(1359) <= "00000000";    
--            LineBuffer0(1360) <= "00000000";
--            LineBuffer0(1361) <= "00000000";
--            LineBuffer0(1362) <= "00000000";
--            LineBuffer0(1363) <= "00000000";
--            LineBuffer0(1364) <= "00000000";
--            LineBuffer0(1365) <= "00000000";
--            LineBuffer0(1366) <= "00000000";
--            LineBuffer0(1367) <= "00000000";
--            LineBuffer0(1368) <= "00000000";
--            LineBuffer0(1369) <= "00000000";    
--            LineBuffer0(1370) <= "00000000";
--            LineBuffer0(1371) <= "00000000";
--            LineBuffer0(1372) <= "00000000";
--            LineBuffer0(1373) <= "00000000";
--            LineBuffer0(1374) <= "00000000";
--            LineBuffer0(1375) <= "00000000";
--            LineBuffer0(1376) <= "00000000";
--            LineBuffer0(1377) <= "00000000";
--            LineBuffer0(1378) <= "00000000";
--            LineBuffer0(1379) <= "00000000";    
--            LineBuffer0(1380) <= "00000000";
--            LineBuffer0(1381) <= "00000000";
--            LineBuffer0(1382) <= "00000000";
--            LineBuffer0(1383) <= "00000000";
--            LineBuffer0(1384) <= "00000000";
--            LineBuffer0(1385) <= "00000000";
--            LineBuffer0(1386) <= "00000000";
--            LineBuffer0(1387) <= "00000000";
--            LineBuffer0(1388) <= "00000000";
--            LineBuffer0(1389) <= "00000000";    
--            LineBuffer0(1390) <= "00000000";
--            LineBuffer0(1391) <= "00000000";
--            LineBuffer0(1392) <= "00000000";
--            LineBuffer0(1393) <= "00000000";
--            LineBuffer0(1394) <= "00000000";
--            LineBuffer0(1395) <= "00000000";
--            LineBuffer0(1396) <= "00000000";
--            LineBuffer0(1397) <= "00000000";
--            LineBuffer0(1398) <= "00000000";
--            LineBuffer0(1399) <= "00000000";    
--            LineBuffer0(1400) <= "00000000";
--            LineBuffer0(1401) <= "00000000";
--            LineBuffer0(1402) <= "00000000";
--            LineBuffer0(1403) <= "00000000";
--            LineBuffer0(1404) <= "00000000";
--            LineBuffer0(1405) <= "00000000";
--            LineBuffer0(1406) <= "00000000";
--            LineBuffer0(1407) <= "00000000";
--            LineBuffer0(1408) <= "00000000";
--            LineBuffer0(1409) <= "00000000";    
--            LineBuffer0(1410) <= "00000000";
--            LineBuffer0(1411) <= "00000000";
--            LineBuffer0(1412) <= "00000000";
--            LineBuffer0(1413) <= "00000000";
--            LineBuffer0(1414) <= "00000000";
--            LineBuffer0(1415) <= "00000000";
--            LineBuffer0(1416) <= "00000000";
--            LineBuffer0(1417) <= "00000000";
--            LineBuffer0(1418) <= "00000000";
--            LineBuffer0(1419) <= "00000000";    
--            LineBuffer0(1420) <= "00000000";
--            LineBuffer0(1421) <= "00000000";
--            LineBuffer0(1422) <= "00000000";
--            LineBuffer0(1423) <= "00000000";
--            LineBuffer0(1424) <= "00000000";
--            LineBuffer0(1425) <= "00000000";
--            LineBuffer0(1426) <= "00000000";
--            LineBuffer0(1427) <= "00000000";
--            LineBuffer0(1428) <= "00000000";
--            LineBuffer0(1429) <= "00000000";    
--            LineBuffer0(1430) <= "00000000";
--            LineBuffer0(1431) <= "00000000";
--            LineBuffer0(1432) <= "00000000";
--            LineBuffer0(1433) <= "00000000";
--            LineBuffer0(1434) <= "00000000";
--            LineBuffer0(1435) <= "00000000";
--            LineBuffer0(1436) <= "00000000";
--            LineBuffer0(1437) <= "00000000";
--            LineBuffer0(1438) <= "00000000";
--            LineBuffer0(1439) <= "00000000";    
--            LineBuffer0(1440) <= "00000000";
--            LineBuffer0(1441) <= "00000000";
--            LineBuffer0(1442) <= "00000000";
--            LineBuffer0(1443) <= "00000000";
--            LineBuffer0(1444) <= "00000000";
--            LineBuffer0(1445) <= "00000000";
--            LineBuffer0(1446) <= "00000000";
--            LineBuffer0(1447) <= "00000000";
--            LineBuffer0(1448) <= "00000000";
--            LineBuffer0(1449) <= "00000000";    
--            LineBuffer0(1450) <= "00000000";
--            LineBuffer0(1451) <= "00000000";
--            LineBuffer0(1452) <= "00000000";
--            LineBuffer0(1453) <= "00000000";
--            LineBuffer0(1454) <= "00000000";
--            LineBuffer0(1455) <= "00000000";
--            LineBuffer0(1456) <= "00000000";
--            LineBuffer0(1457) <= "00000000";
--            LineBuffer0(1458) <= "00000000";
--            LineBuffer0(1459) <= "00000000";    
--            LineBuffer0(1460) <= "00000000";
--            LineBuffer0(1461) <= "00000000";
--            LineBuffer0(1462) <= "00000000";
--            LineBuffer0(1463) <= "00000000";
--            LineBuffer0(1464) <= "00000000";
--            LineBuffer0(1465) <= "00000000";
--            LineBuffer0(1466) <= "00000000";
--            LineBuffer0(1467) <= "00000000";
--            LineBuffer0(1468) <= "00000000";
--            LineBuffer0(1469) <= "00000000";    
--            LineBuffer0(1470) <= "00000000";
--            LineBuffer0(1471) <= "00000000";
--            LineBuffer0(1472) <= "00000000";
--            LineBuffer0(1473) <= "00000000";
--            LineBuffer0(1474) <= "00000000";
--            LineBuffer0(1475) <= "00000000";
--            LineBuffer0(1476) <= "00000000";
--            LineBuffer0(1477) <= "00000000";
--            LineBuffer0(1478) <= "00000000";
--            LineBuffer0(1479) <= "00000000";
--            LineBuffer0(1480) <= "00000000";
--            LineBuffer0(1481) <= "00000000";
--            LineBuffer0(1482) <= "00000000";
--            LineBuffer0(1483) <= "00000000";
--            LineBuffer0(1484) <= "00000000";
--            LineBuffer0(1485) <= "00000000";
--            LineBuffer0(1486) <= "00000000";
--            LineBuffer0(1487) <= "00000000";
--            LineBuffer0(1488) <= "00000000";
--            LineBuffer0(1489) <= "00000000";    
--            LineBuffer0(1490) <= "00000000";
--            LineBuffer0(1491) <= "00000000";
--            LineBuffer0(1492) <= "00000000";
--            LineBuffer0(1493) <= "00000000";
--            LineBuffer0(1494) <= "00000000";
--            LineBuffer0(1495) <= "00000000";
--            LineBuffer0(1496) <= "00000000";
--            LineBuffer0(1497) <= "00000000";
--            LineBuffer0(1498) <= "00000000";
--            LineBuffer0(1499) <= "00000000";    
--            LineBuffer0(1500) <= "00000000";
--            LineBuffer0(1501) <= "00000000";
--            LineBuffer0(1502) <= "00000000";
--            LineBuffer0(1503) <= "00000000";
--            LineBuffer0(1504) <= "00000000";
--            LineBuffer0(1505) <= "00000000";
--            LineBuffer0(1506) <= "00000000";
--            LineBuffer0(1507) <= "00000000";
--            LineBuffer0(1508) <= "00000000";
--            LineBuffer0(1509) <= "00000000";    
--            LineBuffer0(1510) <= "00000000";
--            LineBuffer0(1511) <= "00000000";
--            LineBuffer0(1512) <= "00000000";
--            LineBuffer0(1513) <= "00000000";
--            LineBuffer0(1514) <= "00000000";
--            LineBuffer0(1515) <= "00000000";
--            LineBuffer0(1516) <= "00000000";
--            LineBuffer0(1517) <= "00000000";
--            LineBuffer0(1518) <= "00000000";
--            LineBuffer0(1519) <= "00000000";    
--            LineBuffer0(1520) <= "00000000";
--            LineBuffer0(1521) <= "00000000";
--            LineBuffer0(1522) <= "00000000";
--            LineBuffer0(1523) <= "00000000";
--            LineBuffer0(1524) <= "00000000";
--            LineBuffer0(1525) <= "00000000";
--            LineBuffer0(1526) <= "00000000";
--            LineBuffer0(1527) <= "00000000";
--            LineBuffer0(1528) <= "00000000";
--            LineBuffer0(1529) <= "00000000";    
--            LineBuffer0(1530) <= "00000000";
--            LineBuffer0(1531) <= "00000000";
--            LineBuffer0(1532) <= "00000000";
--            LineBuffer0(1533) <= "00000000";
--            LineBuffer0(1534) <= "00000000";
--            LineBuffer0(1535) <= "00000000";
--            LineBuffer0(1536) <= "00000000";
--            LineBuffer0(1537) <= "00000000";
--            LineBuffer0(1538) <= "00000000";
--            LineBuffer0(1539) <= "00000000";    
--            LineBuffer0(1540) <= "00000000";
--            LineBuffer0(1541) <= "00000000";
--            LineBuffer0(1542) <= "00000000";
--            LineBuffer0(1543) <= "00000000";
--            LineBuffer0(1544) <= "00000000";
--            LineBuffer0(1545) <= "00000000";
--            LineBuffer0(1546) <= "00000000";
--            LineBuffer0(1547) <= "00000000";
--            LineBuffer0(1548) <= "00000000";
--            LineBuffer0(1549) <= "00000000";    
--            LineBuffer0(1550) <= "00000000";
--            LineBuffer0(1551) <= "00000000";
--            LineBuffer0(1552) <= "00000000";
--            LineBuffer0(1553) <= "00000000";
--            LineBuffer0(1554) <= "00000000";
--            LineBuffer0(1555) <= "00000000";
--            LineBuffer0(1556) <= "00000000";
--            LineBuffer0(1557) <= "00000000";
--            LineBuffer0(1558) <= "00000000";
--            LineBuffer0(1559) <= "00000000";    
--            LineBuffer0(1560) <= "00000000";
--            LineBuffer0(1561) <= "00000000";
--            LineBuffer0(1562) <= "00000000";
--            LineBuffer0(1563) <= "00000000";
--            LineBuffer0(1564) <= "00000000";
--            LineBuffer0(1565) <= "00000000";
--            LineBuffer0(1566) <= "00000000";
--            LineBuffer0(1567) <= "00000000";
--            LineBuffer0(1568) <= "00000000";
--            LineBuffer0(1569) <= "00000000";    
--            LineBuffer0(1570) <= "00000000";
--            LineBuffer0(1571) <= "00000000";
--            LineBuffer0(1572) <= "00000000";
--            LineBuffer0(1573) <= "00000000";
--            LineBuffer0(1574) <= "00000000";
--            LineBuffer0(1575) <= "00000000";
--            LineBuffer0(1576) <= "00000000";
--            LineBuffer0(1577) <= "00000000";
--            LineBuffer0(1578) <= "00000000";
--            LineBuffer0(1579) <= "00000000";
--            LineBuffer0(1580) <= "00000000";
--            LineBuffer0(1581) <= "00000000";
--            LineBuffer0(1582) <= "00000000";
--            LineBuffer0(1583) <= "00000000";
--            LineBuffer0(1584) <= "00000000";
--            LineBuffer0(1585) <= "00000000";
--            LineBuffer0(1586) <= "00000000";
--            LineBuffer0(1587) <= "00000000";
--            LineBuffer0(1588) <= "00000000";
--            LineBuffer0(1589) <= "00000000";    
--            LineBuffer0(1590) <= "00000000";
--            LineBuffer0(1591) <= "00000000";
--            LineBuffer0(1592) <= "00000000";
--            LineBuffer0(1593) <= "00000000";
--            LineBuffer0(1594) <= "00000000";
--            LineBuffer0(1595) <= "00000000";
--            LineBuffer0(1596) <= "00000000";
--            LineBuffer0(1597) <= "00000000";
--            LineBuffer0(1598) <= "00000000";
--            LineBuffer0(1599) <= "00000000";    
--            LineBuffer0(1600) <= "00000000";
--            LineBuffer0(1601) <= "00000000";
--            LineBuffer0(1602) <= "00000000";
--            LineBuffer0(1603) <= "00000000";
--            LineBuffer0(1604) <= "00000000";
--            LineBuffer0(1605) <= "00000000";
--            LineBuffer0(1606) <= "00000000";
--            LineBuffer0(1607) <= "00000000";
--            LineBuffer0(1608) <= "00000000";
--            LineBuffer0(1609) <= "00000000";    
--            LineBuffer0(1610) <= "00000000";
--            LineBuffer0(1611) <= "00000000";
--            LineBuffer0(1612) <= "00000000";
--            LineBuffer0(1613) <= "00000000";
--            LineBuffer0(1614) <= "00000000";
--            LineBuffer0(1615) <= "00000000";
--            LineBuffer0(1616) <= "00000000";
--            LineBuffer0(1617) <= "00000000";
--            LineBuffer0(1618) <= "00000000";
--            LineBuffer0(1619) <= "00000000";    
--            LineBuffer0(1620) <= "00000000";
--            LineBuffer0(1621) <= "00000000";
--            LineBuffer0(1622) <= "00000000";
--            LineBuffer0(1623) <= "00000000";
--            LineBuffer0(1624) <= "00000000";
--            LineBuffer0(1625) <= "00000000";
--            LineBuffer0(1626) <= "00000000";
--            LineBuffer0(1627) <= "00000000";
--            LineBuffer0(1628) <= "00000000";
--            LineBuffer0(1629) <= "00000000";    
--            LineBuffer0(1630) <= "00000000";
--            LineBuffer0(1631) <= "00000000";
--            LineBuffer0(1632) <= "00000000";
--            LineBuffer0(1633) <= "00000000";
--            LineBuffer0(1634) <= "00000000";
--            LineBuffer0(1635) <= "00000000";
--            LineBuffer0(1636) <= "00000000";
--            LineBuffer0(1637) <= "00000000";
--            LineBuffer0(1638) <= "00000000";
--            LineBuffer0(1639) <= "00000000";    
--            LineBuffer0(1640) <= "00000000";
--            LineBuffer0(1641) <= "00000000";
--            LineBuffer0(1642) <= "00000000";
--            LineBuffer0(1643) <= "00000000";
--            LineBuffer0(1644) <= "00000000";
--            LineBuffer0(1645) <= "00000000";
--            LineBuffer0(1646) <= "00000000";
--            LineBuffer0(1647) <= "00000000";
--            LineBuffer0(1648) <= "00000000";
--            LineBuffer0(1649) <= "00000000";    
--            LineBuffer0(1650) <= "00000000";
--            LineBuffer0(1651) <= "00000000";
--            LineBuffer0(1652) <= "00000000";
--            LineBuffer0(1653) <= "00000000";
--            LineBuffer0(1654) <= "00000000";
--            LineBuffer0(1655) <= "00000000";
--            LineBuffer0(1656) <= "00000000";
--            LineBuffer0(1657) <= "00000000";
--            LineBuffer0(1658) <= "00000000";
--            LineBuffer0(1659) <= "00000000";    
--            LineBuffer0(1660) <= "00000000";
--            LineBuffer0(1661) <= "00000000";
--            LineBuffer0(1662) <= "00000000";
--            LineBuffer0(1663) <= "00000000";
--            LineBuffer0(1664) <= "00000000";
--            LineBuffer0(1665) <= "00000000";
--            LineBuffer0(1666) <= "00000000";
--            LineBuffer0(1667) <= "00000000";
--            LineBuffer0(1668) <= "00000000";
--            LineBuffer0(1669) <= "00000000";    
--            LineBuffer0(1670) <= "00000000";
--            LineBuffer0(1671) <= "00000000";
--            LineBuffer0(1672) <= "00000000";
--            LineBuffer0(1673) <= "00000000";
--            LineBuffer0(1674) <= "00000000";
--            LineBuffer0(1675) <= "00000000";
--            LineBuffer0(1676) <= "00000000";
--            LineBuffer0(1677) <= "00000000";
--            LineBuffer0(1678) <= "00000000";
--            LineBuffer0(1679) <= "00000000";
--            LineBuffer0(1680) <= "00000000";
--            LineBuffer0(1681) <= "00000000";
--            LineBuffer0(1682) <= "00000000";
--            LineBuffer0(1683) <= "00000000";
--            LineBuffer0(1684) <= "00000000";
--            LineBuffer0(1685) <= "00000000";
--            LineBuffer0(1686) <= "00000000";
--            LineBuffer0(1687) <= "00000000";
--            LineBuffer0(1688) <= "00000000";
--            LineBuffer0(1689) <= "00000000";    
--            LineBuffer0(1690) <= "00000000";
--            LineBuffer0(1691) <= "00000000";
--            LineBuffer0(1692) <= "00000000";
--            LineBuffer0(1693) <= "00000000";
--            LineBuffer0(1694) <= "00000000";
--            LineBuffer0(1695) <= "00000000";
--            LineBuffer0(1696) <= "00000000";
--            LineBuffer0(1697) <= "00000000";
--            LineBuffer0(1698) <= "00000000";
--            LineBuffer0(1699) <= "00000000";    
--            LineBuffer0(1700) <= "00000000";
--            LineBuffer0(1701) <= "00000000";
--            LineBuffer0(1702) <= "00000000";
--            LineBuffer0(1703) <= "00000000";
--            LineBuffer0(1704) <= "00000000";
--            LineBuffer0(1705) <= "00000000";
--            LineBuffer0(1706) <= "00000000";
--            LineBuffer0(1707) <= "00000000";
--            LineBuffer0(1708) <= "00000000";
--            LineBuffer0(1709) <= "00000000";    
--            LineBuffer0(1710) <= "00000000";
--            LineBuffer0(1711) <= "00000000";
--            LineBuffer0(1712) <= "00000000";
--            LineBuffer0(1713) <= "00000000";
--            LineBuffer0(1714) <= "00000000";
--            LineBuffer0(1715) <= "00000000";
--            LineBuffer0(1716) <= "00000000";
--            LineBuffer0(1717) <= "00000000";
--            LineBuffer0(1718) <= "00000000";
--            LineBuffer0(1719) <= "00000000";    
--            LineBuffer0(1720) <= "00000000";
--            LineBuffer0(1721) <= "00000000";
--            LineBuffer0(1722) <= "00000000";
--            LineBuffer0(1723) <= "00000000";
--            LineBuffer0(1724) <= "00000000";
--            LineBuffer0(1725) <= "00000000";
--            LineBuffer0(1726) <= "00000000";
--            LineBuffer0(1727) <= "00000000";
--            LineBuffer0(1728) <= "00000000";
--            LineBuffer0(1729) <= "00000000";    
--            LineBuffer0(1730) <= "00000000";
--            LineBuffer0(1731) <= "00000000";
--            LineBuffer0(1732) <= "00000000";
--            LineBuffer0(1733) <= "00000000";
--            LineBuffer0(1734) <= "00000000";
--            LineBuffer0(1735) <= "00000000";
--            LineBuffer0(1736) <= "00000000";
--            LineBuffer0(1737) <= "00000000";
--            LineBuffer0(1738) <= "00000000";
--            LineBuffer0(1739) <= "00000000";    
--            LineBuffer0(1740) <= "00000000";
--            LineBuffer0(1741) <= "00000000";
--            LineBuffer0(1742) <= "00000000";
--            LineBuffer0(1743) <= "00000000";
--            LineBuffer0(1744) <= "00000000";
--            LineBuffer0(1745) <= "00000000";
--            LineBuffer0(1746) <= "00000000";
--            LineBuffer0(1747) <= "00000000";
--            LineBuffer0(1748) <= "00000000";
--            LineBuffer0(1749) <= "00000000";    
--            LineBuffer0(1750) <= "00000000";
--            LineBuffer0(1751) <= "00000000";
--            LineBuffer0(1752) <= "00000000";
--            LineBuffer0(1753) <= "00000000";
--            LineBuffer0(1754) <= "00000000";
--            LineBuffer0(1755) <= "00000000";
--            LineBuffer0(1756) <= "00000000";
--            LineBuffer0(1757) <= "00000000";
--            LineBuffer0(1758) <= "00000000";
--            LineBuffer0(1759) <= "00000000";    
--            LineBuffer0(1760) <= "00000000";
--            LineBuffer0(1761) <= "00000000";
--            LineBuffer0(1762) <= "00000000";
--            LineBuffer0(1763) <= "00000000";
--            LineBuffer0(1764) <= "00000000";
--            LineBuffer0(1765) <= "00000000";
--            LineBuffer0(1766) <= "00000000";
--            LineBuffer0(1767) <= "00000000";
--            LineBuffer0(1768) <= "00000000";
--            LineBuffer0(1769) <= "00000000";    
--            LineBuffer0(1770) <= "00000000";
--            LineBuffer0(1771) <= "00000000";
--            LineBuffer0(1772) <= "00000000";
--            LineBuffer0(1773) <= "00000000";
--            LineBuffer0(1774) <= "00000000";
--            LineBuffer0(1775) <= "00000000";
--            LineBuffer0(1776) <= "00000000";
--            LineBuffer0(1777) <= "00000000";
--            LineBuffer0(1778) <= "00000000";
--            LineBuffer0(1779) <= "00000000";
--            LineBuffer0(1780) <= "00000000";
--            LineBuffer0(1781) <= "00000000";
--            LineBuffer0(1782) <= "00000000";
--            LineBuffer0(1783) <= "00000000";
--            LineBuffer0(1784) <= "00000000";
--            LineBuffer0(1785) <= "00000000";
--            LineBuffer0(1786) <= "00000000";
--            LineBuffer0(1787) <= "00000000";
--            LineBuffer0(1788) <= "00000000";
--            LineBuffer0(1789) <= "00000000";    
--            LineBuffer0(1790) <= "00000000";
--            LineBuffer0(1791) <= "00000000";
--            LineBuffer0(1792) <= "00000000";
--            LineBuffer0(1793) <= "00000000";
--            LineBuffer0(1794) <= "00000000";
--            LineBuffer0(1795) <= "00000000";
--            LineBuffer0(1796) <= "00000000";
--            LineBuffer0(1797) <= "00000000";
--            LineBuffer0(1798) <= "00000000";
--            LineBuffer0(1799) <= "00000000";    
--            LineBuffer0(1800) <= "00000000";
--            LineBuffer0(1801) <= "00000000";
--            LineBuffer0(1802) <= "00000000";
--            LineBuffer0(1803) <= "00000000";
--            LineBuffer0(1804) <= "00000000";
--            LineBuffer0(1805) <= "00000000";
--            LineBuffer0(1806) <= "00000000";
--            LineBuffer0(1807) <= "00000000";
--            LineBuffer0(1808) <= "00000000";
--            LineBuffer0(1809) <= "00000000";    
--            LineBuffer0(1810) <= "00000000";
--            LineBuffer0(1811) <= "00000000";
--            LineBuffer0(1812) <= "00000000";
--            LineBuffer0(1813) <= "00000000";
--            LineBuffer0(1814) <= "00000000";
--            LineBuffer0(1815) <= "00000000";
--            LineBuffer0(1816) <= "00000000";
--            LineBuffer0(1817) <= "00000000";
--            LineBuffer0(1818) <= "00000000";
--            LineBuffer0(1819) <= "00000000";    
--            LineBuffer0(1820) <= "00000000";
--            LineBuffer0(1821) <= "00000000";
--            LineBuffer0(1822) <= "00000000";
--            LineBuffer0(1823) <= "00000000";
--            LineBuffer0(1824) <= "00000000";
--            LineBuffer0(1825) <= "00000000";
--            LineBuffer0(1826) <= "00000000";
--            LineBuffer0(1827) <= "00000000";
--            LineBuffer0(1828) <= "00000000";
--            LineBuffer0(1829) <= "00000000";    
--            LineBuffer0(1830) <= "00000000";
--            LineBuffer0(1831) <= "00000000";
--            LineBuffer0(1832) <= "00000000";
--            LineBuffer0(1833) <= "00000000";
--            LineBuffer0(1834) <= "00000000";
--            LineBuffer0(1835) <= "00000000";
--            LineBuffer0(1836) <= "00000000";
--            LineBuffer0(1837) <= "00000000";
--            LineBuffer0(1838) <= "00000000";
--            LineBuffer0(1839) <= "00000000";    
--            LineBuffer0(1840) <= "00000000";
--            LineBuffer0(1841) <= "00000000";
--            LineBuffer0(1842) <= "00000000";
--            LineBuffer0(1843) <= "00000000";
--            LineBuffer0(1844) <= "00000000";
--            LineBuffer0(1845) <= "00000000";
--            LineBuffer0(1846) <= "00000000";
--            LineBuffer0(1847) <= "00000000";
--            LineBuffer0(1848) <= "00000000";
--            LineBuffer0(1849) <= "00000000";    
--            LineBuffer0(1850) <= "00000000";
--            LineBuffer0(1851) <= "00000000";
--            LineBuffer0(1852) <= "00000000";
--            LineBuffer0(1853) <= "00000000";
--            LineBuffer0(1854) <= "00000000";
--            LineBuffer0(1855) <= "00000000";
--            LineBuffer0(1856) <= "00000000";
--            LineBuffer0(1857) <= "00000000";
--            LineBuffer0(1858) <= "00000000";
--            LineBuffer0(1859) <= "00000000";    
--            LineBuffer0(1860) <= "00000000";
--            LineBuffer0(1861) <= "00000000";
--            LineBuffer0(1862) <= "00000000";
--            LineBuffer0(1863) <= "00000000";
--            LineBuffer0(1864) <= "00000000";
--            LineBuffer0(1865) <= "00000000";
--            LineBuffer0(1866) <= "00000000";
--            LineBuffer0(1867) <= "00000000";
--            LineBuffer0(1868) <= "00000000";
--            LineBuffer0(1869) <= "00000000";    
--            LineBuffer0(1870) <= "00000000";
--            LineBuffer0(1871) <= "00000000";
--            LineBuffer0(1872) <= "00000000";
--            LineBuffer0(1873) <= "00000000";
--            LineBuffer0(1874) <= "00000000";
--            LineBuffer0(1875) <= "00000000";
--            LineBuffer0(1876) <= "00000000";
--            LineBuffer0(1877) <= "00000000";
--            LineBuffer0(1878) <= "00000000";
--            LineBuffer0(1879) <= "00000000";
--            LineBuffer0(1880) <= "00000000";
--            LineBuffer0(1881) <= "00000000";
--            LineBuffer0(1882) <= "00000000";
--            LineBuffer0(1883) <= "00000000";
--            LineBuffer0(1884) <= "00000000";
--            LineBuffer0(1885) <= "00000000";
--            LineBuffer0(1886) <= "00000000";
--            LineBuffer0(1887) <= "00000000";
--            LineBuffer0(1888) <= "00000000";
--            LineBuffer0(1889) <= "00000000";    
--            LineBuffer0(1890) <= "00000000";
--            LineBuffer0(1891) <= "00000000";
--            LineBuffer0(1892) <= "00000000";
--            LineBuffer0(1893) <= "00000000";
--            LineBuffer0(1894) <= "00000000";
--            LineBuffer0(1895) <= "00000000";
--            LineBuffer0(1896) <= "00000000";
--            LineBuffer0(1897) <= "00000000";
--            LineBuffer0(1898) <= "00000000";
--            LineBuffer0(1899) <= "00000000";    
--            LineBuffer0(1900) <= "00000000";
--            LineBuffer0(1901) <= "00000000";
--            LineBuffer0(1902) <= "00000000";
--            LineBuffer0(1903) <= "00000000";
--            LineBuffer0(1904) <= "00000000";
--            LineBuffer0(1905) <= "00000000";
--            LineBuffer0(1906) <= "00000000";
--            LineBuffer0(1907) <= "00000000";
--            LineBuffer0(1908) <= "00000000";
--            LineBuffer0(1909) <= "00000000";    
--            LineBuffer0(1910) <= "00000000";
--            LineBuffer0(1911) <= "00000000";
--            LineBuffer0(1912) <= "00000000";
--            LineBuffer0(1913) <= "00000000";
--            LineBuffer0(1914) <= "00000000";
--            LineBuffer0(1915) <= "00000000";
--            LineBuffer0(1916) <= "00000000";
--            LineBuffer0(1917) <= "00000000";
--            LineBuffer0(1918) <= "00000000";
--            LineBuffer0(1919) <= "00000000";




		
LineBuffer1(0) <= "00000000";
			LineBuffer1(1) <= "00000000";
			LineBuffer1(2) <= "00000000";
			LineBuffer1(3) <= "00000000";
			LineBuffer1(4) <= "00000000";
			LineBuffer1(5) <= "00000000";
			LineBuffer1(6) <= "00000000";
			LineBuffer1(7) <= "00000000";
			LineBuffer1(8) <= "00000000";
			LineBuffer1(9) <= "00000000";	
			LineBuffer1(10) <= "00000000";
			LineBuffer1(11) <= "00000000";
			LineBuffer1(12) <= "00000000";
			LineBuffer1(13) <= "00000000";
			LineBuffer1(14) <= "00000000";
			LineBuffer1(15) <= "00000000";
			LineBuffer1(16) <= "00000000";
			LineBuffer1(17) <= "00000000";
			LineBuffer1(18) <= "00000000";
			LineBuffer1(19) <= "00000000";	
			LineBuffer1(20) <= "00000000";
			LineBuffer1(21) <= "00000000";
			LineBuffer1(22) <= "00000000";
			LineBuffer1(23) <= "00000000";
			LineBuffer1(24) <= "00000000";
			LineBuffer1(25) <= "00000000";
			LineBuffer1(26) <= "00000000";
			LineBuffer1(27) <= "00000000";
			LineBuffer1(28) <= "00000000";
			LineBuffer1(29) <= "00000000";	
			LineBuffer1(30) <= "00000000";
			LineBuffer1(31) <= "00000000";
			LineBuffer1(32) <= "00000000";
			LineBuffer1(33) <= "00000000";
			LineBuffer1(34) <= "00000000";
			LineBuffer1(35) <= "00000000";
			LineBuffer1(36) <= "00000000";
			LineBuffer1(37) <= "00000000";
			LineBuffer1(38) <= "00000000";
			LineBuffer1(39) <= "00000000";	
			LineBuffer1(40) <= "00000000";
			LineBuffer1(41) <= "00000000";
			LineBuffer1(42) <= "00000000";
			LineBuffer1(43) <= "00000000";
			LineBuffer1(44) <= "00000000";
			LineBuffer1(45) <= "00000000";
			LineBuffer1(46) <= "00000000";
			LineBuffer1(47) <= "00000000";
			LineBuffer1(48) <= "00000000";
			LineBuffer1(49) <= "00000000";	
			LineBuffer1(50) <= "00000000";
			LineBuffer1(51) <= "00000000";
			LineBuffer1(52) <= "00000000";
			LineBuffer1(53) <= "00000000";
			LineBuffer1(54) <= "00000000";
			LineBuffer1(55) <= "00000000";
			LineBuffer1(56) <= "00000000";
			LineBuffer1(57) <= "00000000";
			LineBuffer1(58) <= "00000000";
			LineBuffer1(59) <= "00000000";	
			LineBuffer1(60) <= "00000000";
			LineBuffer1(61) <= "00000000";
			LineBuffer1(62) <= "00000000";
			LineBuffer1(63) <= "00000000";
			LineBuffer1(64) <= "00000000";
			LineBuffer1(65) <= "00000000";
			LineBuffer1(66) <= "00000000";
			LineBuffer1(67) <= "00000000";
			LineBuffer1(68) <= "00000000";
			LineBuffer1(69) <= "00000000";	
			LineBuffer1(70) <= "00000000";
			LineBuffer1(71) <= "00000000";
			LineBuffer1(72) <= "00000000";
			LineBuffer1(73) <= "00000000";
			LineBuffer1(74) <= "00000000";
			LineBuffer1(75) <= "00000000";
			LineBuffer1(76) <= "00000000";
			LineBuffer1(77) <= "00000000";
			LineBuffer1(78) <= "00000000";
			LineBuffer1(79) <= "00000000";	
			LineBuffer1(80) <= "00000000";
			LineBuffer1(81) <= "00000000";
			LineBuffer1(82) <= "00000000";
			LineBuffer1(83) <= "00000000";
			LineBuffer1(84) <= "00000000";
			LineBuffer1(85) <= "00000000";
			LineBuffer1(86) <= "00000000";
			LineBuffer1(87) <= "00000000";
			LineBuffer1(88) <= "00000000";
			LineBuffer1(89) <= "00000000";	
			LineBuffer1(90) <= "00000000";
			LineBuffer1(91) <= "00000000";
			LineBuffer1(92) <= "00000000";
			LineBuffer1(93) <= "00000000";
			LineBuffer1(94) <= "00000000";
			LineBuffer1(95) <= "00000000";
			LineBuffer1(96) <= "00000000";
			LineBuffer1(97) <= "00000000";
			LineBuffer1(98) <= "00000000";
			LineBuffer1(99) <= "00000000";	
			LineBuffer1(100) <= "00000000";
			LineBuffer1(101) <= "00000000";
			LineBuffer1(102) <= "00000000";
			LineBuffer1(103) <= "00000000";
			LineBuffer1(104) <= "00000000";
			LineBuffer1(105) <= "00000000";
			LineBuffer1(106) <= "00000000";
			LineBuffer1(107) <= "00000000";
			LineBuffer1(108) <= "00000000";
			LineBuffer1(109) <= "00000000";	
			LineBuffer1(110) <= "00000000";
			LineBuffer1(111) <= "00000000";
			LineBuffer1(112) <= "00000000";
			LineBuffer1(113) <= "00000000";
			LineBuffer1(114) <= "00000000";
			LineBuffer1(115) <= "00000000";
			LineBuffer1(116) <= "00000000";
			LineBuffer1(117) <= "00000000";
			LineBuffer1(118) <= "00000000";
			LineBuffer1(119) <= "00000000";	
			LineBuffer1(120) <= "00000000";
			LineBuffer1(121) <= "00000000";
			LineBuffer1(122) <= "00000000";
			LineBuffer1(123) <= "00000000";
			LineBuffer1(124) <= "00000000";
			LineBuffer1(125) <= "00000000";
			LineBuffer1(126) <= "00000000";
			LineBuffer1(127) <= "00000000";
			LineBuffer1(128) <= "00000000";
			LineBuffer1(129) <= "00000000";	
			LineBuffer1(130) <= "00000000";
			LineBuffer1(131) <= "00000000";
			LineBuffer1(132) <= "00000000";
			LineBuffer1(133) <= "00000000";
			LineBuffer1(134) <= "00000000";
			LineBuffer1(135) <= "00000000";
			LineBuffer1(136) <= "00000000";
			LineBuffer1(137) <= "00000000";
			LineBuffer1(138) <= "00000000";
			LineBuffer1(139) <= "00000000";	
			LineBuffer1(140) <= "00000000";
			LineBuffer1(141) <= "00000000";
			LineBuffer1(142) <= "00000000";
			LineBuffer1(143) <= "00000000";
			LineBuffer1(144) <= "00000000";
			LineBuffer1(145) <= "00000000";
			LineBuffer1(146) <= "00000000";
			LineBuffer1(147) <= "00000000";
			LineBuffer1(148) <= "00000000";
			LineBuffer1(149) <= "00000000";	
			LineBuffer1(150) <= "00000000";
			LineBuffer1(151) <= "00000000";
			LineBuffer1(152) <= "00000000";
			LineBuffer1(153) <= "00000000";
			LineBuffer1(154) <= "00000000";
			LineBuffer1(155) <= "00000000";
			LineBuffer1(156) <= "00000000";
			LineBuffer1(157) <= "00000000";
			LineBuffer1(158) <= "00000000";
			LineBuffer1(159) <= "00000000";	
			LineBuffer1(160) <= "00000000";
			LineBuffer1(161) <= "00000000";
			LineBuffer1(162) <= "00000000";
			LineBuffer1(163) <= "00000000";
			LineBuffer1(164) <= "00000000";
			LineBuffer1(165) <= "00000000";
			LineBuffer1(166) <= "00000000";
			LineBuffer1(167) <= "00000000";
			LineBuffer1(168) <= "00000000";
			LineBuffer1(169) <= "00000000";	
			LineBuffer1(170) <= "00000000";
			LineBuffer1(171) <= "00000000";
			LineBuffer1(172) <= "00000000";
			LineBuffer1(173) <= "00000000";
			LineBuffer1(174) <= "00000000";
			LineBuffer1(175) <= "00000000";
			LineBuffer1(176) <= "00000000";
			LineBuffer1(177) <= "00000000";
			LineBuffer1(178) <= "00000000";
			LineBuffer1(179) <= "00000000";	
			LineBuffer1(180) <= "00000000";
			LineBuffer1(181) <= "00000000";
			LineBuffer1(182) <= "00000000";
			LineBuffer1(183) <= "00000000";
			LineBuffer1(184) <= "00000000";
			LineBuffer1(185) <= "00000000";
			LineBuffer1(186) <= "00000000";
			LineBuffer1(187) <= "00000000";
			LineBuffer1(188) <= "00000000";
			LineBuffer1(189) <= "00000000";	
			LineBuffer1(190) <= "00000000";
			LineBuffer1(191) <= "00000000";
			LineBuffer1(192) <= "00000000";
			LineBuffer1(193) <= "00000000";
			LineBuffer1(194) <= "00000000";
			LineBuffer1(195) <= "00000000";
			LineBuffer1(196) <= "00000000";
			LineBuffer1(197) <= "00000000";
			LineBuffer1(198) <= "00000000";
			LineBuffer1(199) <= "00000000";
			LineBuffer1(200) <= "00000000";
			LineBuffer1(201) <= "00000000";
			LineBuffer1(202) <= "00000000";
			LineBuffer1(203) <= "00000000";
			LineBuffer1(204) <= "00000000";
			LineBuffer1(205) <= "00000000";
			LineBuffer1(206) <= "00000000";
			LineBuffer1(207) <= "00000000";
			LineBuffer1(208) <= "00000000";
			LineBuffer1(209) <= "00000000";	
			LineBuffer1(210) <= "00000000";
			LineBuffer1(211) <= "00000000";
			LineBuffer1(212) <= "00000000";
			LineBuffer1(213) <= "00000000";
			LineBuffer1(214) <= "00000000";
			LineBuffer1(215) <= "00000000";
			LineBuffer1(216) <= "00000000";
			LineBuffer1(217) <= "00000000";
			LineBuffer1(218) <= "00000000";
			LineBuffer1(219) <= "00000000";	
			LineBuffer1(220) <= "00000000";
			LineBuffer1(221) <= "00000000";
			LineBuffer1(222) <= "00000000";
			LineBuffer1(223) <= "00000000";
			LineBuffer1(224) <= "00000000";
			LineBuffer1(225) <= "00000000";
			LineBuffer1(226) <= "00000000";
			LineBuffer1(227) <= "00000000";
			LineBuffer1(228) <= "00000000";
			LineBuffer1(229) <= "00000000";	
			LineBuffer1(230) <= "00000000";
			LineBuffer1(231) <= "00000000";
			LineBuffer1(232) <= "00000000";
			LineBuffer1(233) <= "00000000";
			LineBuffer1(234) <= "00000000";
			LineBuffer1(235) <= "00000000";
			LineBuffer1(236) <= "00000000";
			LineBuffer1(237) <= "00000000";
			LineBuffer1(238) <= "00000000";
			LineBuffer1(239) <= "00000000";	
			LineBuffer1(240) <= "00000000";
			LineBuffer1(241) <= "00000000";
			LineBuffer1(242) <= "00000000";
			LineBuffer1(243) <= "00000000";
			LineBuffer1(244) <= "00000000";
			LineBuffer1(245) <= "00000000";
			LineBuffer1(246) <= "00000000";
			LineBuffer1(247) <= "00000000";
			LineBuffer1(248) <= "00000000";
			LineBuffer1(249) <= "00000000";	
			LineBuffer1(250) <= "00000000";
			LineBuffer1(251) <= "00000000";
			LineBuffer1(252) <= "00000000";
			LineBuffer1(253) <= "00000000";
			LineBuffer1(254) <= "00000000";
			LineBuffer1(255) <= "00000000";
			LineBuffer1(256) <= "00000000";
			LineBuffer1(257) <= "00000000";
			LineBuffer1(258) <= "00000000";
			LineBuffer1(259) <= "00000000";	
			LineBuffer1(260) <= "00000000";
			LineBuffer1(261) <= "00000000";
			LineBuffer1(262) <= "00000000";
			LineBuffer1(263) <= "00000000";
			LineBuffer1(264) <= "00000000";
			LineBuffer1(265) <= "00000000";
			LineBuffer1(266) <= "00000000";
			LineBuffer1(267) <= "00000000";
			LineBuffer1(268) <= "00000000";
			LineBuffer1(269) <= "00000000";	
			LineBuffer1(270) <= "00000000";
			LineBuffer1(271) <= "00000000";
			LineBuffer1(272) <= "00000000";
			LineBuffer1(273) <= "00000000";
			LineBuffer1(274) <= "00000000";
			LineBuffer1(275) <= "00000000";
			LineBuffer1(276) <= "00000000";
			LineBuffer1(277) <= "00000000";
			LineBuffer1(278) <= "00000000";
			LineBuffer1(279) <= "00000000";	
			LineBuffer1(280) <= "00000000";
			LineBuffer1(281) <= "00000000";
			LineBuffer1(282) <= "00000000";
			LineBuffer1(283) <= "00000000";
			LineBuffer1(284) <= "00000000";
			LineBuffer1(285) <= "00000000";
			LineBuffer1(286) <= "00000000";
			LineBuffer1(287) <= "00000000";
			LineBuffer1(288) <= "00000000";
			LineBuffer1(289) <= "00000000";	
			LineBuffer1(290) <= "00000000";
			LineBuffer1(291) <= "00000000";
			LineBuffer1(292) <= "00000000";
			LineBuffer1(293) <= "00000000";
			LineBuffer1(294) <= "00000000";
			LineBuffer1(295) <= "00000000";
			LineBuffer1(296) <= "00000000";
			LineBuffer1(297) <= "00000000";
			LineBuffer1(298) <= "00000000";
			LineBuffer1(299) <= "00000000";
			LineBuffer1(300) <= "00000000";
			LineBuffer1(301) <= "00000000";
			LineBuffer1(302) <= "00000000";
			LineBuffer1(303) <= "00000000";
			LineBuffer1(304) <= "00000000";
			LineBuffer1(305) <= "00000000";
			LineBuffer1(306) <= "00000000";
			LineBuffer1(307) <= "00000000";
			LineBuffer1(308) <= "00000000";
			LineBuffer1(309) <= "00000000";	
			LineBuffer1(310) <= "00000000";
			LineBuffer1(311) <= "00000000";
			LineBuffer1(312) <= "00000000";
			LineBuffer1(313) <= "00000000";
			LineBuffer1(314) <= "00000000";
			LineBuffer1(315) <= "00000000";
			LineBuffer1(316) <= "00000000";
			LineBuffer1(317) <= "00000000";
			LineBuffer1(318) <= "00000000";
			LineBuffer1(319) <= "00000000";	
			LineBuffer1(320) <= "00000000";
			LineBuffer1(321) <= "00000000";
			LineBuffer1(322) <= "00000000";
			LineBuffer1(323) <= "00000000";
			LineBuffer1(324) <= "00000000";
			LineBuffer1(325) <= "00000000";
			LineBuffer1(326) <= "00000000";
			LineBuffer1(327) <= "00000000";
			LineBuffer1(328) <= "00000000";
			LineBuffer1(329) <= "00000000";	
			LineBuffer1(330) <= "00000000";
			LineBuffer1(331) <= "00000000";
			LineBuffer1(332) <= "00000000";
			LineBuffer1(333) <= "00000000";
			LineBuffer1(334) <= "00000000";
			LineBuffer1(335) <= "00000000";
			LineBuffer1(336) <= "00000000";
			LineBuffer1(337) <= "00000000";
			LineBuffer1(338) <= "00000000";
			LineBuffer1(339) <= "00000000";	
			LineBuffer1(340) <= "00000000";
			LineBuffer1(341) <= "00000000";
			LineBuffer1(342) <= "00000000";
			LineBuffer1(343) <= "00000000";
			LineBuffer1(344) <= "00000000";
			LineBuffer1(345) <= "00000000";
			LineBuffer1(346) <= "00000000";
			LineBuffer1(347) <= "00000000";
			LineBuffer1(348) <= "00000000";
			LineBuffer1(349) <= "00000000";	
			LineBuffer1(350) <= "00000000";
			LineBuffer1(351) <= "00000000";
			LineBuffer1(352) <= "00000000";
			LineBuffer1(353) <= "00000000";
			LineBuffer1(354) <= "00000000";
			LineBuffer1(355) <= "00000000";
			LineBuffer1(356) <= "00000000";
			LineBuffer1(357) <= "00000000";
			LineBuffer1(358) <= "00000000";
			LineBuffer1(359) <= "00000000";	
			LineBuffer1(360) <= "00000000";
			LineBuffer1(361) <= "00000000";
			LineBuffer1(362) <= "00000000";
			LineBuffer1(363) <= "00000000";
			LineBuffer1(364) <= "00000000";
			LineBuffer1(365) <= "00000000";
			LineBuffer1(366) <= "00000000";
			LineBuffer1(367) <= "00000000";
			LineBuffer1(368) <= "00000000";
			LineBuffer1(369) <= "00000000";	
			LineBuffer1(370) <= "00000000";
			LineBuffer1(371) <= "00000000";
			LineBuffer1(372) <= "00000000";
			LineBuffer1(373) <= "00000000";
			LineBuffer1(374) <= "00000000";
			LineBuffer1(375) <= "00000000";
			LineBuffer1(376) <= "00000000";
			LineBuffer1(377) <= "00000000";
			LineBuffer1(378) <= "00000000";
			LineBuffer1(379) <= "00000000";	
			LineBuffer1(380) <= "00000000";
			LineBuffer1(381) <= "00000000";
			LineBuffer1(382) <= "00000000";
			LineBuffer1(383) <= "00000000";
			LineBuffer1(384) <= "00000000";
			LineBuffer1(385) <= "00000000";
			LineBuffer1(386) <= "00000000";
			LineBuffer1(387) <= "00000000";
			LineBuffer1(388) <= "00000000";
			LineBuffer1(389) <= "00000000";	
			LineBuffer1(390) <= "00000000";
			LineBuffer1(391) <= "00000000";
			LineBuffer1(392) <= "00000000";
			LineBuffer1(393) <= "00000000";
			LineBuffer1(394) <= "00000000";
			LineBuffer1(395) <= "00000000";
			LineBuffer1(396) <= "00000000";
			LineBuffer1(397) <= "00000000";
			LineBuffer1(398) <= "00000000";
			LineBuffer1(399) <= "00000000";
			LineBuffer1(400) <= "00000000";
			LineBuffer1(401) <= "00000000";
			LineBuffer1(402) <= "00000000";
			LineBuffer1(403) <= "00000000";
			LineBuffer1(404) <= "00000000";
			LineBuffer1(405) <= "00000000";
			LineBuffer1(406) <= "00000000";
			LineBuffer1(407) <= "00000000";
			LineBuffer1(408) <= "00000000";
			LineBuffer1(409) <= "00000000";	
			LineBuffer1(410) <= "00000000";
			LineBuffer1(411) <= "00000000";
			LineBuffer1(412) <= "00000000";
			LineBuffer1(413) <= "00000000";
			LineBuffer1(414) <= "00000000";
			LineBuffer1(415) <= "00000000";
			LineBuffer1(416) <= "00000000";
			LineBuffer1(417) <= "00000000";
			LineBuffer1(418) <= "00000000";
			LineBuffer1(419) <= "00000000";	
			LineBuffer1(420) <= "00000000";
			LineBuffer1(421) <= "00000000";
			LineBuffer1(422) <= "00000000";
			LineBuffer1(423) <= "00000000";
			LineBuffer1(424) <= "00000000";
			LineBuffer1(425) <= "00000000";
			LineBuffer1(426) <= "00000000";
			LineBuffer1(427) <= "00000000";
			LineBuffer1(428) <= "00000000";
			LineBuffer1(429) <= "00000000";	
			LineBuffer1(430) <= "00000000";
			LineBuffer1(431) <= "00000000";
			LineBuffer1(432) <= "00000000";
			LineBuffer1(433) <= "00000000";
			LineBuffer1(434) <= "00000000";
			LineBuffer1(435) <= "00000000";
			LineBuffer1(436) <= "00000000";
			LineBuffer1(437) <= "00000000";
			LineBuffer1(438) <= "00000000";
			LineBuffer1(439) <= "00000000";	
			LineBuffer1(440) <= "00000000";
			LineBuffer1(441) <= "00000000";
			LineBuffer1(442) <= "00000000";
			LineBuffer1(443) <= "00000000";
			LineBuffer1(444) <= "00000000";
			LineBuffer1(445) <= "00000000";
			LineBuffer1(446) <= "00000000";
			LineBuffer1(447) <= "00000000";
			LineBuffer1(448) <= "00000000";
			LineBuffer1(449) <= "00000000";	
			LineBuffer1(450) <= "00000000";
			LineBuffer1(451) <= "00000000";
			LineBuffer1(452) <= "00000000";
			LineBuffer1(453) <= "00000000";
			LineBuffer1(454) <= "00000000";
			LineBuffer1(455) <= "00000000";
			LineBuffer1(456) <= "00000000";
			LineBuffer1(457) <= "00000000";
			LineBuffer1(458) <= "00000000";
			LineBuffer1(459) <= "00000000";	
			LineBuffer1(460) <= "00000000";
			LineBuffer1(461) <= "00000000";
			LineBuffer1(462) <= "00000000";
			LineBuffer1(463) <= "00000000";
			LineBuffer1(464) <= "00000000";
			LineBuffer1(465) <= "00000000";
			LineBuffer1(466) <= "00000000";
			LineBuffer1(467) <= "00000000";
			LineBuffer1(468) <= "00000000";
			LineBuffer1(469) <= "00000000";	
			LineBuffer1(470) <= "00000000";
			LineBuffer1(471) <= "00000000";
			LineBuffer1(472) <= "00000000";
			LineBuffer1(473) <= "00000000";
			LineBuffer1(474) <= "00000000";
			LineBuffer1(475) <= "00000000";
			LineBuffer1(476) <= "00000000";
			LineBuffer1(477) <= "00000000";
			LineBuffer1(478) <= "00000000";
			LineBuffer1(479) <= "00000000";	
			LineBuffer1(480) <= "00000000";
			LineBuffer1(481) <= "00000000";
			LineBuffer1(482) <= "00000000";
			LineBuffer1(483) <= "00000000";
			LineBuffer1(484) <= "00000000";
			LineBuffer1(485) <= "00000000";
			LineBuffer1(486) <= "00000000";
			LineBuffer1(487) <= "00000000";
			LineBuffer1(488) <= "00000000";
			LineBuffer1(489) <= "00000000";	
			LineBuffer1(490) <= "00000000";
			LineBuffer1(491) <= "00000000";
			LineBuffer1(492) <= "00000000";
			LineBuffer1(493) <= "00000000";
			LineBuffer1(494) <= "00000000";
			LineBuffer1(495) <= "00000000";
			LineBuffer1(496) <= "00000000";
			LineBuffer1(497) <= "00000000";
			LineBuffer1(498) <= "00000000";
			LineBuffer1(499) <= "00000000";
			LineBuffer1(500) <= "00000000";
			LineBuffer1(501) <= "00000000";
			LineBuffer1(502) <= "00000000";
			LineBuffer1(503) <= "00000000";
			LineBuffer1(504) <= "00000000";
			LineBuffer1(505) <= "00000000";
			LineBuffer1(506) <= "00000000";
			LineBuffer1(507) <= "00000000";
			LineBuffer1(508) <= "00000000";
			LineBuffer1(509) <= "00000000";	
			LineBuffer1(510) <= "00000000";
			LineBuffer1(511) <= "00000000";
			LineBuffer1(512) <= "00000000";
			LineBuffer1(513) <= "00000000";
			LineBuffer1(514) <= "00000000";
			LineBuffer1(515) <= "00000000";
			LineBuffer1(516) <= "00000000";
			LineBuffer1(517) <= "00000000";
			LineBuffer1(518) <= "00000000";
			LineBuffer1(519) <= "00000000";	
			LineBuffer1(520) <= "00000000";
			LineBuffer1(521) <= "00000000";
			LineBuffer1(522) <= "00000000";
			LineBuffer1(523) <= "00000000";
			LineBuffer1(524) <= "00000000";
			LineBuffer1(525) <= "00000000";
			LineBuffer1(526) <= "00000000";
			LineBuffer1(527) <= "00000000";
			LineBuffer1(528) <= "00000000";
			LineBuffer1(529) <= "00000000";	
			LineBuffer1(530) <= "00000000";
			LineBuffer1(531) <= "00000000";
			LineBuffer1(532) <= "00000000";
			LineBuffer1(533) <= "00000000";
			LineBuffer1(534) <= "00000000";
			LineBuffer1(535) <= "00000000";
			LineBuffer1(536) <= "00000000";
			LineBuffer1(537) <= "00000000";
			LineBuffer1(538) <= "00000000";
			LineBuffer1(539) <= "00000000";	
			LineBuffer1(540) <= "00000000";
			LineBuffer1(541) <= "00000000";
			LineBuffer1(542) <= "00000000";
			LineBuffer1(543) <= "00000000";
			LineBuffer1(544) <= "00000000";
			LineBuffer1(545) <= "00000000";
			LineBuffer1(546) <= "00000000";
			LineBuffer1(547) <= "00000000";
			LineBuffer1(548) <= "00000000";
			LineBuffer1(549) <= "00000000";	
			LineBuffer1(550) <= "00000000";
			LineBuffer1(551) <= "00000000";
			LineBuffer1(552) <= "00000000";
			LineBuffer1(553) <= "00000000";
			LineBuffer1(554) <= "00000000";
			LineBuffer1(555) <= "00000000";
			LineBuffer1(556) <= "00000000";
			LineBuffer1(557) <= "00000000";
			LineBuffer1(558) <= "00000000";
			LineBuffer1(559) <= "00000000";	
			LineBuffer1(560) <= "00000000";
			LineBuffer1(561) <= "00000000";
			LineBuffer1(562) <= "00000000";
			LineBuffer1(563) <= "00000000";
			LineBuffer1(564) <= "00000000";
			LineBuffer1(565) <= "00000000";
			LineBuffer1(566) <= "00000000";
			LineBuffer1(567) <= "00000000";
			LineBuffer1(568) <= "00000000";
			LineBuffer1(569) <= "00000000";	
			LineBuffer1(570) <= "00000000";
			LineBuffer1(571) <= "00000000";
			LineBuffer1(572) <= "00000000";
			LineBuffer1(573) <= "00000000";
			LineBuffer1(574) <= "00000000";
			LineBuffer1(575) <= "00000000";
			LineBuffer1(576) <= "00000000";
			LineBuffer1(577) <= "00000000";
			LineBuffer1(578) <= "00000000";
			LineBuffer1(579) <= "00000000";	
			LineBuffer1(580) <= "00000000";
			LineBuffer1(581) <= "00000000";
			LineBuffer1(582) <= "00000000";
			LineBuffer1(583) <= "00000000";
			LineBuffer1(584) <= "00000000";
			LineBuffer1(585) <= "00000000";
			LineBuffer1(586) <= "00000000";
			LineBuffer1(587) <= "00000000";
			LineBuffer1(588) <= "00000000";
			LineBuffer1(589) <= "00000000";	
			LineBuffer1(590) <= "00000000";
			LineBuffer1(591) <= "00000000";
			LineBuffer1(592) <= "00000000";
			LineBuffer1(593) <= "00000000";
			LineBuffer1(594) <= "00000000";
			LineBuffer1(595) <= "00000000";
			LineBuffer1(596) <= "00000000";
			LineBuffer1(597) <= "00000000";
			LineBuffer1(598) <= "00000000";
			LineBuffer1(599) <= "00000000";
			LineBuffer1(600) <= "00000000";
			LineBuffer1(601) <= "00000000";
			LineBuffer1(602) <= "00000000";
			LineBuffer1(603) <= "00000000";
			LineBuffer1(604) <= "00000000";
			LineBuffer1(605) <= "00000000";
			LineBuffer1(606) <= "00000000";
			LineBuffer1(607) <= "00000000";
			LineBuffer1(608) <= "00000000";
			LineBuffer1(609) <= "00000000";	
			LineBuffer1(610) <= "00000000";
			LineBuffer1(611) <= "00000000";
			LineBuffer1(612) <= "00000000";
			LineBuffer1(613) <= "00000000";
			LineBuffer1(614) <= "00000000";
			LineBuffer1(615) <= "00000000";
			LineBuffer1(616) <= "00000000";
			LineBuffer1(617) <= "00000000";
			LineBuffer1(618) <= "00000000";
			LineBuffer1(619) <= "00000000";	
			LineBuffer1(620) <= "00000000";
			LineBuffer1(621) <= "00000000";
			LineBuffer1(622) <= "00000000";
			LineBuffer1(623) <= "00000000";
			LineBuffer1(624) <= "00000000";
			LineBuffer1(625) <= "00000000";
			LineBuffer1(626) <= "00000000";
			LineBuffer1(627) <= "00000000";
			LineBuffer1(628) <= "00000000";
			LineBuffer1(629) <= "00000000";	
			LineBuffer1(630) <= "00000000";
			LineBuffer1(631) <= "00000000";
			LineBuffer1(632) <= "00000000";
			LineBuffer1(633) <= "00000000";
			LineBuffer1(634) <= "00000000";
			LineBuffer1(635) <= "00000000";
			LineBuffer1(636) <= "00000000";
			LineBuffer1(637) <= "00000000";
			LineBuffer1(638) <= "00000000";
			LineBuffer1(639) <= "00000000";
			LineBuffer1(640) <= "00000000";
            LineBuffer1(641) <= "00000000";
            LineBuffer1(642) <= "00000000";
            LineBuffer1(643) <= "00000000";
            LineBuffer1(644) <= "00000000";
            LineBuffer1(645) <= "00000000";
            LineBuffer1(646) <= "00000000";
            LineBuffer1(647) <= "00000000";
            LineBuffer1(648) <= "00000000";
            LineBuffer1(649) <= "00000000";    
            LineBuffer1(650) <= "00000000";
            LineBuffer1(651) <= "00000000";
            LineBuffer1(652) <= "00000000";
            LineBuffer1(653) <= "00000000";
            LineBuffer1(654) <= "00000000";
            LineBuffer1(655) <= "00000000";
            LineBuffer1(656) <= "00000000";
            LineBuffer1(657) <= "00000000";
            LineBuffer1(658) <= "00000000";
            LineBuffer1(659) <= "00000000";    
            LineBuffer1(660) <= "00000000";
            LineBuffer1(661) <= "00000000";
            LineBuffer1(662) <= "00000000";
            LineBuffer1(663) <= "00000000";
            LineBuffer1(664) <= "00000000";
            LineBuffer1(665) <= "00000000";
            LineBuffer1(666) <= "00000000";
            LineBuffer1(667) <= "00000000";
            LineBuffer1(668) <= "00000000";
            LineBuffer1(669) <= "00000000";    
            LineBuffer1(670) <= "00000000";
            LineBuffer1(671) <= "00000000";
            LineBuffer1(672) <= "00000000";
            LineBuffer1(673) <= "00000000";
            LineBuffer1(674) <= "00000000";
            LineBuffer1(675) <= "00000000";
            LineBuffer1(676) <= "00000000";
            LineBuffer1(677) <= "00000000";
            LineBuffer1(678) <= "00000000";
            LineBuffer1(679) <= "00000000";    
            LineBuffer1(680) <= "00000000";
            LineBuffer1(681) <= "00000000";
            LineBuffer1(682) <= "00000000";
            LineBuffer1(683) <= "00000000";
            LineBuffer1(684) <= "00000000";
            LineBuffer1(685) <= "00000000";
            LineBuffer1(686) <= "00000000";
            LineBuffer1(687) <= "00000000";
            LineBuffer1(688) <= "00000000";
            LineBuffer1(689) <= "00000000";    
            LineBuffer1(690) <= "00000000";
            LineBuffer1(691) <= "00000000";
            LineBuffer1(692) <= "00000000";
            LineBuffer1(693) <= "00000000";
            LineBuffer1(694) <= "00000000";
            LineBuffer1(695) <= "00000000";
            LineBuffer1(696) <= "00000000";
            LineBuffer1(697) <= "00000000";
            LineBuffer1(698) <= "00000000";
            LineBuffer1(699) <= "00000000";    
            LineBuffer1(700) <= "00000000";
            LineBuffer1(701) <= "00000000";
            LineBuffer1(702) <= "00000000";
            LineBuffer1(703) <= "00000000";
            LineBuffer1(704) <= "00000000";
            LineBuffer1(705) <= "00000000";
            LineBuffer1(706) <= "00000000";
            LineBuffer1(707) <= "00000000";
            LineBuffer1(708) <= "00000000";
            LineBuffer1(709) <= "00000000";    
            LineBuffer1(710) <= "00000000";
            LineBuffer1(711) <= "00000000";
            LineBuffer1(712) <= "00000000";
            LineBuffer1(713) <= "00000000";
            LineBuffer1(714) <= "00000000";
            LineBuffer1(715) <= "00000000";
            LineBuffer1(716) <= "00000000";
            LineBuffer1(717) <= "00000000";
            LineBuffer1(718) <= "00000000";
            LineBuffer1(719) <= "00000000";    
            LineBuffer1(720) <= "00000000";
            LineBuffer1(721) <= "00000000";
            LineBuffer1(722) <= "00000000";
            LineBuffer1(723) <= "00000000";
            LineBuffer1(724) <= "00000000";
            LineBuffer1(725) <= "00000000";
            LineBuffer1(726) <= "00000000";
            LineBuffer1(727) <= "00000000";
            LineBuffer1(728) <= "00000000";
            LineBuffer1(729) <= "00000000";    
            LineBuffer1(730) <= "00000000";
            LineBuffer1(731) <= "00000000";
            LineBuffer1(732) <= "00000000";
            LineBuffer1(733) <= "00000000";
            LineBuffer1(734) <= "00000000";
            LineBuffer1(735) <= "00000000";
            LineBuffer1(736) <= "00000000";
            LineBuffer1(737) <= "00000000";
            LineBuffer1(738) <= "00000000";
            LineBuffer1(739) <= "00000000";    
            LineBuffer1(740) <= "00000000";
            LineBuffer1(741) <= "00000000";
            LineBuffer1(742) <= "00000000";
            LineBuffer1(743) <= "00000000";
            LineBuffer1(744) <= "00000000";
            LineBuffer1(745) <= "00000000";
            LineBuffer1(746) <= "00000000";
            LineBuffer1(747) <= "00000000";
            LineBuffer1(748) <= "00000000";
            LineBuffer1(749) <= "00000000";    
            LineBuffer1(750) <= "00000000";
            LineBuffer1(751) <= "00000000";
            LineBuffer1(752) <= "00000000";
            LineBuffer1(753) <= "00000000";
            LineBuffer1(754) <= "00000000";
            LineBuffer1(755) <= "00000000";
            LineBuffer1(756) <= "00000000";
            LineBuffer1(757) <= "00000000";
            LineBuffer1(758) <= "00000000";
            LineBuffer1(759) <= "00000000";    
            LineBuffer1(760) <= "00000000";
            LineBuffer1(761) <= "00000000";
            LineBuffer1(762) <= "00000000";
            LineBuffer1(763) <= "00000000";
            LineBuffer1(764) <= "00000000";
            LineBuffer1(765) <= "00000000";
            LineBuffer1(766) <= "00000000";
            LineBuffer1(767) <= "00000000";
            LineBuffer1(768) <= "00000000";
            LineBuffer1(769) <= "00000000";    
            LineBuffer1(770) <= "00000000";
            LineBuffer1(771) <= "00000000";
            LineBuffer1(772) <= "00000000";
            LineBuffer1(773) <= "00000000";
            LineBuffer1(774) <= "00000000";
            LineBuffer1(775) <= "00000000";
            LineBuffer1(776) <= "00000000";
            LineBuffer1(777) <= "00000000";
            LineBuffer1(778) <= "00000000";
            LineBuffer1(779) <= "00000000";    
            LineBuffer1(780) <= "00000000";
            LineBuffer1(781) <= "00000000";
            LineBuffer1(782) <= "00000000";
            LineBuffer1(783) <= "00000000";
            LineBuffer1(784) <= "00000000";
            LineBuffer1(785) <= "00000000";
            LineBuffer1(786) <= "00000000";
            LineBuffer1(787) <= "00000000";
            LineBuffer1(788) <= "00000000";
            LineBuffer1(789) <= "00000000";    
            LineBuffer1(790) <= "00000000";
            LineBuffer1(791) <= "00000000";
            LineBuffer1(792) <= "00000000";
            LineBuffer1(793) <= "00000000";
            LineBuffer1(794) <= "00000000";
            LineBuffer1(795) <= "00000000";
            LineBuffer1(796) <= "00000000";
            LineBuffer1(797) <= "00000000";
            LineBuffer1(798) <= "00000000";
            LineBuffer1(799) <= "00000000";    
            LineBuffer1(800) <= "00000000";
            LineBuffer1(801) <= "00000000";
            LineBuffer1(802) <= "00000000";
            LineBuffer1(803) <= "00000000";
            LineBuffer1(804) <= "00000000";
            LineBuffer1(805) <= "00000000";
            LineBuffer1(806) <= "00000000";
            LineBuffer1(807) <= "00000000";
            LineBuffer1(808) <= "00000000";
            LineBuffer1(809) <= "00000000";    
            LineBuffer1(810) <= "00000000";
            LineBuffer1(811) <= "00000000";
            LineBuffer1(812) <= "00000000";
            LineBuffer1(813) <= "00000000";
            LineBuffer1(814) <= "00000000";
            LineBuffer1(815) <= "00000000";
            LineBuffer1(816) <= "00000000";
            LineBuffer1(817) <= "00000000";
            LineBuffer1(818) <= "00000000";
            LineBuffer1(819) <= "00000000";    
            LineBuffer1(820) <= "00000000";
            LineBuffer1(821) <= "00000000";
            LineBuffer1(822) <= "00000000";
            LineBuffer1(823) <= "00000000";
            LineBuffer1(824) <= "00000000";
            LineBuffer1(825) <= "00000000";
            LineBuffer1(826) <= "00000000";
            LineBuffer1(827) <= "00000000";
            LineBuffer1(828) <= "00000000";
            LineBuffer1(829) <= "00000000";    
            LineBuffer1(830) <= "00000000";
            LineBuffer1(831) <= "00000000";
            LineBuffer1(832) <= "00000000";
            LineBuffer1(833) <= "00000000";
            LineBuffer1(834) <= "00000000";
            LineBuffer1(835) <= "00000000";
            LineBuffer1(836) <= "00000000";
            LineBuffer1(837) <= "00000000";
            LineBuffer1(838) <= "00000000";
            LineBuffer1(839) <= "00000000";
            LineBuffer1(840) <= "00000000";
            LineBuffer1(841) <= "00000000";
            LineBuffer1(842) <= "00000000";
            LineBuffer1(843) <= "00000000";
            LineBuffer1(844) <= "00000000";
            LineBuffer1(845) <= "00000000";
            LineBuffer1(846) <= "00000000";
            LineBuffer1(847) <= "00000000";
            LineBuffer1(848) <= "00000000";
            LineBuffer1(849) <= "00000000";    
            LineBuffer1(850) <= "00000000";
            LineBuffer1(851) <= "00000000";
            LineBuffer1(852) <= "00000000";
            LineBuffer1(853) <= "00000000";
            LineBuffer1(854) <= "00000000";
            LineBuffer1(855) <= "00000000";
            LineBuffer1(856) <= "00000000";
            LineBuffer1(857) <= "00000000";
            LineBuffer1(858) <= "00000000";
            LineBuffer1(859) <= "00000000";    
            LineBuffer1(860) <= "00000000";
            LineBuffer1(861) <= "00000000";
            LineBuffer1(862) <= "00000000";
            LineBuffer1(863) <= "00000000";
            LineBuffer1(864) <= "00000000";
            LineBuffer1(865) <= "00000000";
            LineBuffer1(866) <= "00000000";
            LineBuffer1(867) <= "00000000";
            LineBuffer1(868) <= "00000000";
            LineBuffer1(869) <= "00000000";    
            LineBuffer1(870) <= "00000000";
            LineBuffer1(871) <= "00000000";
            LineBuffer1(872) <= "00000000";
            LineBuffer1(873) <= "00000000";
            LineBuffer1(874) <= "00000000";
            LineBuffer1(875) <= "00000000";
            LineBuffer1(876) <= "00000000";
            LineBuffer1(877) <= "00000000";
            LineBuffer1(878) <= "00000000";
            LineBuffer1(879) <= "00000000";    
            LineBuffer1(880) <= "00000000";
            LineBuffer1(881) <= "00000000";
            LineBuffer1(882) <= "00000000";
            LineBuffer1(883) <= "00000000";
            LineBuffer1(884) <= "00000000";
            LineBuffer1(885) <= "00000000";
            LineBuffer1(886) <= "00000000";
            LineBuffer1(887) <= "00000000";
            LineBuffer1(888) <= "00000000";
            LineBuffer1(889) <= "00000000";    
            LineBuffer1(890) <= "00000000";
            LineBuffer1(891) <= "00000000";
            LineBuffer1(892) <= "00000000";
            LineBuffer1(893) <= "00000000";
            LineBuffer1(894) <= "00000000";
            LineBuffer1(895) <= "00000000";
            LineBuffer1(896) <= "00000000";
            LineBuffer1(897) <= "00000000";
            LineBuffer1(898) <= "00000000";
            LineBuffer1(899) <= "00000000";    
            LineBuffer1(900) <= "00000000";
            LineBuffer1(901) <= "00000000";
            LineBuffer1(902) <= "00000000";
            LineBuffer1(903) <= "00000000";
            LineBuffer1(904) <= "00000000";
            LineBuffer1(905) <= "00000000";
            LineBuffer1(906) <= "00000000";
            LineBuffer1(907) <= "00000000";
            LineBuffer1(908) <= "00000000";
            LineBuffer1(909) <= "00000000";    
            LineBuffer1(910) <= "00000000";
            LineBuffer1(911) <= "00000000";
            LineBuffer1(912) <= "00000000";
            LineBuffer1(913) <= "00000000";
            LineBuffer1(914) <= "00000000";
            LineBuffer1(915) <= "00000000";
            LineBuffer1(916) <= "00000000";
            LineBuffer1(917) <= "00000000";
            LineBuffer1(918) <= "00000000";
            LineBuffer1(919) <= "00000000";    
            LineBuffer1(920) <= "00000000";
            LineBuffer1(921) <= "00000000";
            LineBuffer1(922) <= "00000000";
            LineBuffer1(923) <= "00000000";
            LineBuffer1(924) <= "00000000";
            LineBuffer1(925) <= "00000000";
            LineBuffer1(926) <= "00000000";
            LineBuffer1(927) <= "00000000";
            LineBuffer1(928) <= "00000000";
            LineBuffer1(929) <= "00000000";    
            LineBuffer1(930) <= "00000000";
            LineBuffer1(931) <= "00000000";
            LineBuffer1(932) <= "00000000";
            LineBuffer1(933) <= "00000000";
            LineBuffer1(934) <= "00000000";
            LineBuffer1(935) <= "00000000";
            LineBuffer1(936) <= "00000000";
            LineBuffer1(937) <= "00000000";
            LineBuffer1(938) <= "00000000";
            LineBuffer1(939) <= "00000000";
            LineBuffer1(940) <= "00000000";
            LineBuffer1(941) <= "00000000";
            LineBuffer1(942) <= "00000000";
            LineBuffer1(943) <= "00000000";
            LineBuffer1(944) <= "00000000";
            LineBuffer1(945) <= "00000000";
            LineBuffer1(946) <= "00000000";
            LineBuffer1(947) <= "00000000";
            LineBuffer1(948) <= "00000000";
            LineBuffer1(949) <= "00000000";    
            LineBuffer1(950) <= "00000000";
            LineBuffer1(951) <= "00000000";
            LineBuffer1(952) <= "00000000";
            LineBuffer1(953) <= "00000000";
            LineBuffer1(954) <= "00000000";
            LineBuffer1(955) <= "00000000";
            LineBuffer1(956) <= "00000000";
            LineBuffer1(957) <= "00000000";
            LineBuffer1(958) <= "00000000";
            LineBuffer1(959) <= "00000000";    
            LineBuffer1(960) <= "00000000";
            LineBuffer1(961) <= "00000000";
            LineBuffer1(962) <= "00000000";
            LineBuffer1(963) <= "00000000";
            LineBuffer1(964) <= "00000000";
            LineBuffer1(965) <= "00000000";
            LineBuffer1(966) <= "00000000";
            LineBuffer1(967) <= "00000000";
            LineBuffer1(968) <= "00000000";
            LineBuffer1(969) <= "00000000";    
            LineBuffer1(970) <= "00000000";
            LineBuffer1(971) <= "00000000";
            LineBuffer1(972) <= "00000000";
            LineBuffer1(973) <= "00000000";
            LineBuffer1(974) <= "00000000";
            LineBuffer1(975) <= "00000000";
            LineBuffer1(976) <= "00000000";
            LineBuffer1(977) <= "00000000";
            LineBuffer1(978) <= "00000000";
            LineBuffer1(979) <= "00000000";    
            LineBuffer1(980) <= "00000000";
            LineBuffer1(981) <= "00000000";
            LineBuffer1(982) <= "00000000";
            LineBuffer1(983) <= "00000000";
            LineBuffer1(984) <= "00000000";
            LineBuffer1(985) <= "00000000";
            LineBuffer1(986) <= "00000000";
            LineBuffer1(987) <= "00000000";
            LineBuffer1(988) <= "00000000";
            LineBuffer1(989) <= "00000000";    
            LineBuffer1(990) <= "00000000";
            LineBuffer1(991) <= "00000000";
            LineBuffer1(992) <= "00000000";
            LineBuffer1(993) <= "00000000";
            LineBuffer1(994) <= "00000000";
            LineBuffer1(995) <= "00000000";
            LineBuffer1(996) <= "00000000";
            LineBuffer1(997) <= "00000000";
            LineBuffer1(998) <= "00000000";
            LineBuffer1(999) <= "00000000";    
            LineBuffer1(1000) <= "00000000";
            LineBuffer1(1001) <= "00000000";
            LineBuffer1(1002) <= "00000000";
            LineBuffer1(1003) <= "00000000";
            LineBuffer1(1004) <= "00000000";
            LineBuffer1(1005) <= "00000000";
            LineBuffer1(1006) <= "00000000";
            LineBuffer1(1007) <= "00000000";
            LineBuffer1(1008) <= "00000000";
            LineBuffer1(1009) <= "00000000";    
            LineBuffer1(1010) <= "00000000";
            LineBuffer1(1011) <= "00000000";
            LineBuffer1(1012) <= "00000000";
            LineBuffer1(1013) <= "00000000";
            LineBuffer1(1014) <= "00000000";
            LineBuffer1(1015) <= "00000000";
            LineBuffer1(1016) <= "00000000";
            LineBuffer1(1017) <= "00000000";
            LineBuffer1(1018) <= "00000000";
            LineBuffer1(1019) <= "00000000";    
            LineBuffer1(1020) <= "00000000";
            LineBuffer1(1021) <= "00000000";
            LineBuffer1(1022) <= "00000000";
            LineBuffer1(1023) <= "00000000";
            LineBuffer1(1024) <= "00000000";
            LineBuffer1(1025) <= "00000000";
            LineBuffer1(1026) <= "00000000";
            LineBuffer1(1027) <= "00000000";
            LineBuffer1(1028) <= "00000000";
            LineBuffer1(1029) <= "00000000";    
            LineBuffer1(1030) <= "00000000";
            LineBuffer1(1031) <= "00000000";
            LineBuffer1(1032) <= "00000000";
            LineBuffer1(1033) <= "00000000";
            LineBuffer1(1034) <= "00000000";
            LineBuffer1(1035) <= "00000000";
            LineBuffer1(1036) <= "00000000";
            LineBuffer1(1037) <= "00000000";
            LineBuffer1(1038) <= "00000000";
            LineBuffer1(1039) <= "00000000";
            LineBuffer1(1040) <= "00000000";
            LineBuffer1(1041) <= "00000000";
            LineBuffer1(1042) <= "00000000";
            LineBuffer1(1043) <= "00000000";
            LineBuffer1(1044) <= "00000000";
            LineBuffer1(1045) <= "00000000";
            LineBuffer1(1046) <= "00000000";
            LineBuffer1(1047) <= "00000000";
            LineBuffer1(1048) <= "00000000";
            LineBuffer1(1049) <= "00000000";    
            LineBuffer1(1050) <= "00000000";
            LineBuffer1(1051) <= "00000000";
            LineBuffer1(1052) <= "00000000";
            LineBuffer1(1053) <= "00000000";
            LineBuffer1(1054) <= "00000000";
            LineBuffer1(1055) <= "00000000";
            LineBuffer1(1056) <= "00000000";
            LineBuffer1(1057) <= "00000000";
            LineBuffer1(1058) <= "00000000";
            LineBuffer1(1059) <= "00000000";    
            LineBuffer1(1060) <= "00000000";
            LineBuffer1(1061) <= "00000000";
            LineBuffer1(1062) <= "00000000";
            LineBuffer1(1063) <= "00000000";
            LineBuffer1(1064) <= "00000000";
            LineBuffer1(1065) <= "00000000";
            LineBuffer1(1066) <= "00000000";
            LineBuffer1(1067) <= "00000000";
            LineBuffer1(1068) <= "00000000";
            LineBuffer1(1069) <= "00000000";    
            LineBuffer1(1070) <= "00000000";
            LineBuffer1(1071) <= "00000000";
            LineBuffer1(1072) <= "00000000";
            LineBuffer1(1073) <= "00000000";
            LineBuffer1(1074) <= "00000000";
            LineBuffer1(1075) <= "00000000";
            LineBuffer1(1076) <= "00000000";
            LineBuffer1(1077) <= "00000000";
            LineBuffer1(1078) <= "00000000";
            LineBuffer1(1079) <= "00000000";    
            LineBuffer1(1080) <= "00000000";
            LineBuffer1(1081) <= "00000000";
            LineBuffer1(1082) <= "00000000";
            LineBuffer1(1083) <= "00000000";
            LineBuffer1(1084) <= "00000000";
            LineBuffer1(1085) <= "00000000";
            LineBuffer1(1086) <= "00000000";
            LineBuffer1(1087) <= "00000000";
            LineBuffer1(1088) <= "00000000";
            LineBuffer1(1089) <= "00000000";    
            LineBuffer1(1090) <= "00000000";
            LineBuffer1(1091) <= "00000000";
            LineBuffer1(1092) <= "00000000";
            LineBuffer1(1093) <= "00000000";
            LineBuffer1(1094) <= "00000000";
            LineBuffer1(1095) <= "00000000";
            LineBuffer1(1096) <= "00000000";
            LineBuffer1(1097) <= "00000000";
            LineBuffer1(1098) <= "00000000";
            LineBuffer1(1099) <= "00000000";    
            LineBuffer1(1100) <= "00000000";
            LineBuffer1(1101) <= "00000000";
            LineBuffer1(1102) <= "00000000";
            LineBuffer1(1103) <= "00000000";
            LineBuffer1(1104) <= "00000000";
            LineBuffer1(1105) <= "00000000";
            LineBuffer1(1106) <= "00000000";
            LineBuffer1(1107) <= "00000000";
            LineBuffer1(1108) <= "00000000";
            LineBuffer1(1109) <= "00000000";    
            LineBuffer1(1110) <= "00000000";
            LineBuffer1(1111) <= "00000000";
            LineBuffer1(1112) <= "00000000";
            LineBuffer1(1113) <= "00000000";
            LineBuffer1(1114) <= "00000000";
            LineBuffer1(1115) <= "00000000";
            LineBuffer1(1116) <= "00000000";
            LineBuffer1(1117) <= "00000000";
            LineBuffer1(1118) <= "00000000";
            LineBuffer1(1119) <= "00000000";    
            LineBuffer1(1120) <= "00000000";
            LineBuffer1(1121) <= "00000000";
            LineBuffer1(1122) <= "00000000";
            LineBuffer1(1123) <= "00000000";
            LineBuffer1(1124) <= "00000000";
            LineBuffer1(1125) <= "00000000";
            LineBuffer1(1126) <= "00000000";
            LineBuffer1(1127) <= "00000000";
            LineBuffer1(1128) <= "00000000";
            LineBuffer1(1129) <= "00000000";    
            LineBuffer1(1130) <= "00000000";
            LineBuffer1(1131) <= "00000000";
            LineBuffer1(1132) <= "00000000";
            LineBuffer1(1133) <= "00000000";
            LineBuffer1(1134) <= "00000000";
            LineBuffer1(1135) <= "00000000";
            LineBuffer1(1136) <= "00000000";
            LineBuffer1(1137) <= "00000000";
            LineBuffer1(1138) <= "00000000";
            LineBuffer1(1139) <= "00000000";
            LineBuffer1(1140) <= "00000000";
            LineBuffer1(1141) <= "00000000";
            LineBuffer1(1142) <= "00000000";
            LineBuffer1(1143) <= "00000000";
            LineBuffer1(1144) <= "00000000";
            LineBuffer1(1145) <= "00000000";
            LineBuffer1(1146) <= "00000000";
            LineBuffer1(1147) <= "00000000";
            LineBuffer1(1148) <= "00000000";
            LineBuffer1(1149) <= "00000000";    
            LineBuffer1(1150) <= "00000000";
            LineBuffer1(1151) <= "00000000";
            LineBuffer1(1152) <= "00000000";
            LineBuffer1(1153) <= "00000000";
            LineBuffer1(1154) <= "00000000";
            LineBuffer1(1155) <= "00000000";
            LineBuffer1(1156) <= "00000000";
            LineBuffer1(1157) <= "00000000";
            LineBuffer1(1158) <= "00000000";
            LineBuffer1(1159) <= "00000000";    
            LineBuffer1(1160) <= "00000000";
            LineBuffer1(1161) <= "00000000";
            LineBuffer1(1162) <= "00000000";
            LineBuffer1(1163) <= "00000000";
            LineBuffer1(1164) <= "00000000";
            LineBuffer1(1165) <= "00000000";
            LineBuffer1(1166) <= "00000000";
            LineBuffer1(1167) <= "00000000";
            LineBuffer1(1168) <= "00000000";
            LineBuffer1(1169) <= "00000000";    
            LineBuffer1(1170) <= "00000000";
            LineBuffer1(1171) <= "00000000";
            LineBuffer1(1172) <= "00000000";
            LineBuffer1(1173) <= "00000000";
            LineBuffer1(1174) <= "00000000";
            LineBuffer1(1175) <= "00000000";
            LineBuffer1(1176) <= "00000000";
            LineBuffer1(1177) <= "00000000";
            LineBuffer1(1178) <= "00000000";
            LineBuffer1(1179) <= "00000000";    
            LineBuffer1(1180) <= "00000000";
            LineBuffer1(1181) <= "00000000";
            LineBuffer1(1182) <= "00000000";
            LineBuffer1(1183) <= "00000000";
            LineBuffer1(1184) <= "00000000";
            LineBuffer1(1185) <= "00000000";
            LineBuffer1(1186) <= "00000000";
            LineBuffer1(1187) <= "00000000";
            LineBuffer1(1188) <= "00000000";
            LineBuffer1(1189) <= "00000000";    
            LineBuffer1(1190) <= "00000000";
            LineBuffer1(1191) <= "00000000";
            LineBuffer1(1192) <= "00000000";
            LineBuffer1(1193) <= "00000000";
            LineBuffer1(1194) <= "00000000";
            LineBuffer1(1195) <= "00000000";
            LineBuffer1(1196) <= "00000000";
            LineBuffer1(1197) <= "00000000";
            LineBuffer1(1198) <= "00000000";
            LineBuffer1(1199) <= "00000000";    
            LineBuffer1(1200) <= "00000000";
            LineBuffer1(1201) <= "00000000";
            LineBuffer1(1202) <= "00000000";
            LineBuffer1(1203) <= "00000000";
            LineBuffer1(1204) <= "00000000";
            LineBuffer1(1205) <= "00000000";
            LineBuffer1(1206) <= "00000000";
            LineBuffer1(1207) <= "00000000";
            LineBuffer1(1208) <= "00000000";
            LineBuffer1(1209) <= "00000000";    
            LineBuffer1(1210) <= "00000000";
            LineBuffer1(1211) <= "00000000";
            LineBuffer1(1212) <= "00000000";
            LineBuffer1(1213) <= "00000000";
            LineBuffer1(1214) <= "00000000";
            LineBuffer1(1215) <= "00000000";
            LineBuffer1(1216) <= "00000000";
            LineBuffer1(1217) <= "00000000";
            LineBuffer1(1218) <= "00000000";
            LineBuffer1(1219) <= "00000000";    
            LineBuffer1(1220) <= "00000000";
            LineBuffer1(1221) <= "00000000";
            LineBuffer1(1222) <= "00000000";
            LineBuffer1(1223) <= "00000000";
            LineBuffer1(1224) <= "00000000";
            LineBuffer1(1225) <= "00000000";
            LineBuffer1(1226) <= "00000000";
            LineBuffer1(1227) <= "00000000";
            LineBuffer1(1228) <= "00000000";
            LineBuffer1(1229) <= "00000000";    
            LineBuffer1(1230) <= "00000000";
            LineBuffer1(1231) <= "00000000";
            LineBuffer1(1232) <= "00000000";
            LineBuffer1(1233) <= "00000000";
            LineBuffer1(1234) <= "00000000";
            LineBuffer1(1235) <= "00000000";
            LineBuffer1(1236) <= "00000000";
            LineBuffer1(1237) <= "00000000";
            LineBuffer1(1238) <= "00000000";
            LineBuffer1(1239) <= "00000000";
            LineBuffer1(1240) <= "00000000";
            LineBuffer1(1241) <= "00000000";
            LineBuffer1(1242) <= "00000000";
            LineBuffer1(1243) <= "00000000";
            LineBuffer1(1244) <= "00000000";
            LineBuffer1(1245) <= "00000000";
            LineBuffer1(1246) <= "00000000";
            LineBuffer1(1247) <= "00000000";
            LineBuffer1(1248) <= "00000000";
            LineBuffer1(1249) <= "00000000";    
            LineBuffer1(1250) <= "00000000";
            LineBuffer1(1251) <= "00000000";
            LineBuffer1(1252) <= "00000000";
            LineBuffer1(1253) <= "00000000";
            LineBuffer1(1254) <= "00000000";
            LineBuffer1(1255) <= "00000000";
            LineBuffer1(1256) <= "00000000";
            LineBuffer1(1257) <= "00000000";
            LineBuffer1(1258) <= "00000000";
            LineBuffer1(1259) <= "00000000";    
            LineBuffer1(1260) <= "00000000";
            LineBuffer1(1261) <= "00000000";
            LineBuffer1(1262) <= "00000000";
            LineBuffer1(1263) <= "00000000";
            LineBuffer1(1264) <= "00000000";
            LineBuffer1(1265) <= "00000000";
            LineBuffer1(1266) <= "00000000";
            LineBuffer1(1267) <= "00000000";
            LineBuffer1(1268) <= "00000000";
            LineBuffer1(1269) <= "00000000";    
            LineBuffer1(1270) <= "00000000";
            LineBuffer1(1271) <= "00000000";
            LineBuffer1(1272) <= "00000000";
            LineBuffer1(1273) <= "00000000";
            LineBuffer1(1274) <= "00000000";
            LineBuffer1(1275) <= "00000000";
            LineBuffer1(1276) <= "00000000";
            LineBuffer1(1277) <= "00000000";
            LineBuffer1(1278) <= "00000000";
            LineBuffer1(1279) <= "00000000";
            
            
--            LineBuffer1(1280) <= "00000000";
--            LineBuffer1(1281) <= "00000000";
--            LineBuffer1(1282) <= "00000000";
--            LineBuffer1(1283) <= "00000000";
--            LineBuffer1(1284) <= "00000000";
--            LineBuffer1(1285) <= "00000000";
--            LineBuffer1(1286) <= "00000000";
--            LineBuffer1(1287) <= "00000000";
--            LineBuffer1(1288) <= "00000000";
--            LineBuffer1(1289) <= "00000000";    
--            LineBuffer1(1290) <= "00000000";
--            LineBuffer1(1291) <= "00000000";
--            LineBuffer1(1292) <= "00000000";
--            LineBuffer1(1293) <= "00000000";
--            LineBuffer1(1294) <= "00000000";
--            LineBuffer1(1295) <= "00000000";
--            LineBuffer1(1296) <= "00000000";
--            LineBuffer1(1297) <= "00000000";
--            LineBuffer1(1298) <= "00000000";
--            LineBuffer1(1299) <= "00000000";    
--            LineBuffer1(1300) <= "00000000";
--            LineBuffer1(1301) <= "00000000";
--            LineBuffer1(1302) <= "00000000";
--            LineBuffer1(1303) <= "00000000";
--            LineBuffer1(1304) <= "00000000";
--            LineBuffer1(1305) <= "00000000";
--            LineBuffer1(1306) <= "00000000";
--            LineBuffer1(1307) <= "00000000";
--            LineBuffer1(1308) <= "00000000";
--            LineBuffer1(1309) <= "00000000";    
--            LineBuffer1(1310) <= "00000000";
--            LineBuffer1(1311) <= "00000000";
--            LineBuffer1(1312) <= "00000000";
--            LineBuffer1(1313) <= "00000000";
--            LineBuffer1(1314) <= "00000000";
--            LineBuffer1(1315) <= "00000000";
--            LineBuffer1(1316) <= "00000000";
--            LineBuffer1(1317) <= "00000000";
--            LineBuffer1(1318) <= "00000000";
--            LineBuffer1(1319) <= "00000000";    
--            LineBuffer1(1320) <= "00000000";
--            LineBuffer1(1321) <= "00000000";
--            LineBuffer1(1322) <= "00000000";
--            LineBuffer1(1323) <= "00000000";
--            LineBuffer1(1324) <= "00000000";
--            LineBuffer1(1325) <= "00000000";
--            LineBuffer1(1326) <= "00000000";
--            LineBuffer1(1327) <= "00000000";
--            LineBuffer1(1328) <= "00000000";
--            LineBuffer1(1329) <= "00000000";    
--            LineBuffer1(1330) <= "00000000";
--            LineBuffer1(1331) <= "00000000";
--            LineBuffer1(1332) <= "00000000";
--            LineBuffer1(1333) <= "00000000";
--            LineBuffer1(1334) <= "00000000";
--            LineBuffer1(1335) <= "00000000";
--            LineBuffer1(1336) <= "00000000";
--            LineBuffer1(1337) <= "00000000";
--            LineBuffer1(1338) <= "00000000";
--            LineBuffer1(1339) <= "00000000";    
--            LineBuffer1(1340) <= "00000000";
--            LineBuffer1(1341) <= "00000000";
--            LineBuffer1(1342) <= "00000000";
--            LineBuffer1(1343) <= "00000000";
--            LineBuffer1(1344) <= "00000000";
--            LineBuffer1(1345) <= "00000000";
--            LineBuffer1(1346) <= "00000000";
--            LineBuffer1(1347) <= "00000000";
--            LineBuffer1(1348) <= "00000000";
--            LineBuffer1(1349) <= "00000000";    
--            LineBuffer1(1350) <= "00000000";
--            LineBuffer1(1351) <= "00000000";
--            LineBuffer1(1352) <= "00000000";
--            LineBuffer1(1353) <= "00000000";
--            LineBuffer1(1354) <= "00000000";
--            LineBuffer1(1355) <= "00000000";
--            LineBuffer1(1356) <= "00000000";
--            LineBuffer1(1357) <= "00000000";
--            LineBuffer1(1358) <= "00000000";
--            LineBuffer1(1359) <= "00000000";    
--            LineBuffer1(1360) <= "00000000";
--            LineBuffer1(1361) <= "00000000";
--            LineBuffer1(1362) <= "00000000";
--            LineBuffer1(1363) <= "00000000";
--            LineBuffer1(1364) <= "00000000";
--            LineBuffer1(1365) <= "00000000";
--            LineBuffer1(1366) <= "00000000";
--            LineBuffer1(1367) <= "00000000";
--            LineBuffer1(1368) <= "00000000";
--            LineBuffer1(1369) <= "00000000";    
--            LineBuffer1(1370) <= "00000000";
--            LineBuffer1(1371) <= "00000000";
--            LineBuffer1(1372) <= "00000000";
--            LineBuffer1(1373) <= "00000000";
--            LineBuffer1(1374) <= "00000000";
--            LineBuffer1(1375) <= "00000000";
--            LineBuffer1(1376) <= "00000000";
--            LineBuffer1(1377) <= "00000000";
--            LineBuffer1(1378) <= "00000000";
--            LineBuffer1(1379) <= "00000000";    
--            LineBuffer1(1380) <= "00000000";
--            LineBuffer1(1381) <= "00000000";
--            LineBuffer1(1382) <= "00000000";
--            LineBuffer1(1383) <= "00000000";
--            LineBuffer1(1384) <= "00000000";
--            LineBuffer1(1385) <= "00000000";
--            LineBuffer1(1386) <= "00000000";
--            LineBuffer1(1387) <= "00000000";
--            LineBuffer1(1388) <= "00000000";
--            LineBuffer1(1389) <= "00000000";    
--            LineBuffer1(1390) <= "00000000";
--            LineBuffer1(1391) <= "00000000";
--            LineBuffer1(1392) <= "00000000";
--            LineBuffer1(1393) <= "00000000";
--            LineBuffer1(1394) <= "00000000";
--            LineBuffer1(1395) <= "00000000";
--            LineBuffer1(1396) <= "00000000";
--            LineBuffer1(1397) <= "00000000";
--            LineBuffer1(1398) <= "00000000";
--            LineBuffer1(1399) <= "00000000";    
--            LineBuffer1(1400) <= "00000000";
--            LineBuffer1(1401) <= "00000000";
--            LineBuffer1(1402) <= "00000000";
--            LineBuffer1(1403) <= "00000000";
--            LineBuffer1(1404) <= "00000000";
--            LineBuffer1(1405) <= "00000000";
--            LineBuffer1(1406) <= "00000000";
--            LineBuffer1(1407) <= "00000000";
--            LineBuffer1(1408) <= "00000000";
--            LineBuffer1(1409) <= "00000000";    
--            LineBuffer1(1410) <= "00000000";
--            LineBuffer1(1411) <= "00000000";
--            LineBuffer1(1412) <= "00000000";
--            LineBuffer1(1413) <= "00000000";
--            LineBuffer1(1414) <= "00000000";
--            LineBuffer1(1415) <= "00000000";
--            LineBuffer1(1416) <= "00000000";
--            LineBuffer1(1417) <= "00000000";
--            LineBuffer1(1418) <= "00000000";
--            LineBuffer1(1419) <= "00000000";    
--            LineBuffer1(1420) <= "00000000";
--            LineBuffer1(1421) <= "00000000";
--            LineBuffer1(1422) <= "00000000";
--            LineBuffer1(1423) <= "00000000";
--            LineBuffer1(1424) <= "00000000";
--            LineBuffer1(1425) <= "00000000";
--            LineBuffer1(1426) <= "00000000";
--            LineBuffer1(1427) <= "00000000";
--            LineBuffer1(1428) <= "00000000";
--            LineBuffer1(1429) <= "00000000";    
--            LineBuffer1(1430) <= "00000000";
--            LineBuffer1(1431) <= "00000000";
--            LineBuffer1(1432) <= "00000000";
--            LineBuffer1(1433) <= "00000000";
--            LineBuffer1(1434) <= "00000000";
--            LineBuffer1(1435) <= "00000000";
--            LineBuffer1(1436) <= "00000000";
--            LineBuffer1(1437) <= "00000000";
--            LineBuffer1(1438) <= "00000000";
--            LineBuffer1(1439) <= "00000000";    
--            LineBuffer1(1440) <= "00000000";
--            LineBuffer1(1441) <= "00000000";
--            LineBuffer1(1442) <= "00000000";
--            LineBuffer1(1443) <= "00000000";
--            LineBuffer1(1444) <= "00000000";
--            LineBuffer1(1445) <= "00000000";
--            LineBuffer1(1446) <= "00000000";
--            LineBuffer1(1447) <= "00000000";
--            LineBuffer1(1448) <= "00000000";
--            LineBuffer1(1449) <= "00000000";    
--            LineBuffer1(1450) <= "00000000";
--            LineBuffer1(1451) <= "00000000";
--            LineBuffer1(1452) <= "00000000";
--            LineBuffer1(1453) <= "00000000";
--            LineBuffer1(1454) <= "00000000";
--            LineBuffer1(1455) <= "00000000";
--            LineBuffer1(1456) <= "00000000";
--            LineBuffer1(1457) <= "00000000";
--            LineBuffer1(1458) <= "00000000";
--            LineBuffer1(1459) <= "00000000";    
--            LineBuffer1(1460) <= "00000000";
--            LineBuffer1(1461) <= "00000000";
--            LineBuffer1(1462) <= "00000000";
--            LineBuffer1(1463) <= "00000000";
--            LineBuffer1(1464) <= "00000000";
--            LineBuffer1(1465) <= "00000000";
--            LineBuffer1(1466) <= "00000000";
--            LineBuffer1(1467) <= "00000000";
--            LineBuffer1(1468) <= "00000000";
--            LineBuffer1(1469) <= "00000000";    
--            LineBuffer1(1470) <= "00000000";
--            LineBuffer1(1471) <= "00000000";
--            LineBuffer1(1472) <= "00000000";
--            LineBuffer1(1473) <= "00000000";
--            LineBuffer1(1474) <= "00000000";
--            LineBuffer1(1475) <= "00000000";
--            LineBuffer1(1476) <= "00000000";
--            LineBuffer1(1477) <= "00000000";
--            LineBuffer1(1478) <= "00000000";
--            LineBuffer1(1479) <= "00000000";
--            LineBuffer1(1480) <= "00000000";
--            LineBuffer1(1481) <= "00000000";
--            LineBuffer1(1482) <= "00000000";
--            LineBuffer1(1483) <= "00000000";
--            LineBuffer1(1484) <= "00000000";
--            LineBuffer1(1485) <= "00000000";
--            LineBuffer1(1486) <= "00000000";
--            LineBuffer1(1487) <= "00000000";
--            LineBuffer1(1488) <= "00000000";
--            LineBuffer1(1489) <= "00000000";    
--            LineBuffer1(1490) <= "00000000";
--            LineBuffer1(1491) <= "00000000";
--            LineBuffer1(1492) <= "00000000";
--            LineBuffer1(1493) <= "00000000";
--            LineBuffer1(1494) <= "00000000";
--            LineBuffer1(1495) <= "00000000";
--            LineBuffer1(1496) <= "00000000";
--            LineBuffer1(1497) <= "00000000";
--            LineBuffer1(1498) <= "00000000";
--            LineBuffer1(1499) <= "00000000";    
--            LineBuffer1(1500) <= "00000000";
--            LineBuffer1(1501) <= "00000000";
--            LineBuffer1(1502) <= "00000000";
--            LineBuffer1(1503) <= "00000000";
--            LineBuffer1(1504) <= "00000000";
--            LineBuffer1(1505) <= "00000000";
--            LineBuffer1(1506) <= "00000000";
--            LineBuffer1(1507) <= "00000000";
--            LineBuffer1(1508) <= "00000000";
--            LineBuffer1(1509) <= "00000000";    
--            LineBuffer1(1510) <= "00000000";
--            LineBuffer1(1511) <= "00000000";
--            LineBuffer1(1512) <= "00000000";
--            LineBuffer1(1513) <= "00000000";
--            LineBuffer1(1514) <= "00000000";
--            LineBuffer1(1515) <= "00000000";
--            LineBuffer1(1516) <= "00000000";
--            LineBuffer1(1517) <= "00000000";
--            LineBuffer1(1518) <= "00000000";
--            LineBuffer1(1519) <= "00000000";    
--            LineBuffer1(1520) <= "00000000";
--            LineBuffer1(1521) <= "00000000";
--            LineBuffer1(1522) <= "00000000";
--            LineBuffer1(1523) <= "00000000";
--            LineBuffer1(1524) <= "00000000";
--            LineBuffer1(1525) <= "00000000";
--            LineBuffer1(1526) <= "00000000";
--            LineBuffer1(1527) <= "00000000";
--            LineBuffer1(1528) <= "00000000";
--            LineBuffer1(1529) <= "00000000";    
--            LineBuffer1(1530) <= "00000000";
--            LineBuffer1(1531) <= "00000000";
--            LineBuffer1(1532) <= "00000000";
--            LineBuffer1(1533) <= "00000000";
--            LineBuffer1(1534) <= "00000000";
--            LineBuffer1(1535) <= "00000000";
--            LineBuffer1(1536) <= "00000000";
--            LineBuffer1(1537) <= "00000000";
--            LineBuffer1(1538) <= "00000000";
--            LineBuffer1(1539) <= "00000000";    
--            LineBuffer1(1540) <= "00000000";
--            LineBuffer1(1541) <= "00000000";
--            LineBuffer1(1542) <= "00000000";
--            LineBuffer1(1543) <= "00000000";
--            LineBuffer1(1544) <= "00000000";
--            LineBuffer1(1545) <= "00000000";
--            LineBuffer1(1546) <= "00000000";
--            LineBuffer1(1547) <= "00000000";
--            LineBuffer1(1548) <= "00000000";
--            LineBuffer1(1549) <= "00000000";    
--            LineBuffer1(1550) <= "00000000";
--            LineBuffer1(1551) <= "00000000";
--            LineBuffer1(1552) <= "00000000";
--            LineBuffer1(1553) <= "00000000";
--            LineBuffer1(1554) <= "00000000";
--            LineBuffer1(1555) <= "00000000";
--            LineBuffer1(1556) <= "00000000";
--            LineBuffer1(1557) <= "00000000";
--            LineBuffer1(1558) <= "00000000";
--            LineBuffer1(1559) <= "00000000";    
--            LineBuffer1(1560) <= "00000000";
--            LineBuffer1(1561) <= "00000000";
--            LineBuffer1(1562) <= "00000000";
--            LineBuffer1(1563) <= "00000000";
--            LineBuffer1(1564) <= "00000000";
--            LineBuffer1(1565) <= "00000000";
--            LineBuffer1(1566) <= "00000000";
--            LineBuffer1(1567) <= "00000000";
--            LineBuffer1(1568) <= "00000000";
--            LineBuffer1(1569) <= "00000000";    
--            LineBuffer1(1570) <= "00000000";
--            LineBuffer1(1571) <= "00000000";
--            LineBuffer1(1572) <= "00000000";
--            LineBuffer1(1573) <= "00000000";
--            LineBuffer1(1574) <= "00000000";
--            LineBuffer1(1575) <= "00000000";
--            LineBuffer1(1576) <= "00000000";
--            LineBuffer1(1577) <= "00000000";
--            LineBuffer1(1578) <= "00000000";
--            LineBuffer1(1579) <= "00000000";
--            LineBuffer1(1580) <= "00000000";
--            LineBuffer1(1581) <= "00000000";
--            LineBuffer1(1582) <= "00000000";
--            LineBuffer1(1583) <= "00000000";
--            LineBuffer1(1584) <= "00000000";
--            LineBuffer1(1585) <= "00000000";
--            LineBuffer1(1586) <= "00000000";
--            LineBuffer1(1587) <= "00000000";
--            LineBuffer1(1588) <= "00000000";
--            LineBuffer1(1589) <= "00000000";    
--            LineBuffer1(1590) <= "00000000";
--            LineBuffer1(1591) <= "00000000";
--            LineBuffer1(1592) <= "00000000";
--            LineBuffer1(1593) <= "00000000";
--            LineBuffer1(1594) <= "00000000";
--            LineBuffer1(1595) <= "00000000";
--            LineBuffer1(1596) <= "00000000";
--            LineBuffer1(1597) <= "00000000";
--            LineBuffer1(1598) <= "00000000";
--            LineBuffer1(1599) <= "00000000";    
--            LineBuffer1(1600) <= "00000000";
--            LineBuffer1(1601) <= "00000000";
--            LineBuffer1(1602) <= "00000000";
--            LineBuffer1(1603) <= "00000000";
--            LineBuffer1(1604) <= "00000000";
--            LineBuffer1(1605) <= "00000000";
--            LineBuffer1(1606) <= "00000000";
--            LineBuffer1(1607) <= "00000000";
--            LineBuffer1(1608) <= "00000000";
--            LineBuffer1(1609) <= "00000000";    
--            LineBuffer1(1610) <= "00000000";
--            LineBuffer1(1611) <= "00000000";
--            LineBuffer1(1612) <= "00000000";
--            LineBuffer1(1613) <= "00000000";
--            LineBuffer1(1614) <= "00000000";
--            LineBuffer1(1615) <= "00000000";
--            LineBuffer1(1616) <= "00000000";
--            LineBuffer1(1617) <= "00000000";
--            LineBuffer1(1618) <= "00000000";
--            LineBuffer1(1619) <= "00000000";    
--            LineBuffer1(1620) <= "00000000";
--            LineBuffer1(1621) <= "00000000";
--            LineBuffer1(1622) <= "00000000";
--            LineBuffer1(1623) <= "00000000";
--            LineBuffer1(1624) <= "00000000";
--            LineBuffer1(1625) <= "00000000";
--            LineBuffer1(1626) <= "00000000";
--            LineBuffer1(1627) <= "00000000";
--            LineBuffer1(1628) <= "00000000";
--            LineBuffer1(1629) <= "00000000";    
--            LineBuffer1(1630) <= "00000000";
--            LineBuffer1(1631) <= "00000000";
--            LineBuffer1(1632) <= "00000000";
--            LineBuffer1(1633) <= "00000000";
--            LineBuffer1(1634) <= "00000000";
--            LineBuffer1(1635) <= "00000000";
--            LineBuffer1(1636) <= "00000000";
--            LineBuffer1(1637) <= "00000000";
--            LineBuffer1(1638) <= "00000000";
--            LineBuffer1(1639) <= "00000000";    
--            LineBuffer1(1640) <= "00000000";
--            LineBuffer1(1641) <= "00000000";
--            LineBuffer1(1642) <= "00000000";
--            LineBuffer1(1643) <= "00000000";
--            LineBuffer1(1644) <= "00000000";
--            LineBuffer1(1645) <= "00000000";
--            LineBuffer1(1646) <= "00000000";
--            LineBuffer1(1647) <= "00000000";
--            LineBuffer1(1648) <= "00000000";
--            LineBuffer1(1649) <= "00000000";    
--            LineBuffer1(1650) <= "00000000";
--            LineBuffer1(1651) <= "00000000";
--            LineBuffer1(1652) <= "00000000";
--            LineBuffer1(1653) <= "00000000";
--            LineBuffer1(1654) <= "00000000";
--            LineBuffer1(1655) <= "00000000";
--            LineBuffer1(1656) <= "00000000";
--            LineBuffer1(1657) <= "00000000";
--            LineBuffer1(1658) <= "00000000";
--            LineBuffer1(1659) <= "00000000";    
--            LineBuffer1(1660) <= "00000000";
--            LineBuffer1(1661) <= "00000000";
--            LineBuffer1(1662) <= "00000000";
--            LineBuffer1(1663) <= "00000000";
--            LineBuffer1(1664) <= "00000000";
--            LineBuffer1(1665) <= "00000000";
--            LineBuffer1(1666) <= "00000000";
--            LineBuffer1(1667) <= "00000000";
--            LineBuffer1(1668) <= "00000000";
--            LineBuffer1(1669) <= "00000000";    
--            LineBuffer1(1670) <= "00000000";
--            LineBuffer1(1671) <= "00000000";
--            LineBuffer1(1672) <= "00000000";
--            LineBuffer1(1673) <= "00000000";
--            LineBuffer1(1674) <= "00000000";
--            LineBuffer1(1675) <= "00000000";
--            LineBuffer1(1676) <= "00000000";
--            LineBuffer1(1677) <= "00000000";
--            LineBuffer1(1678) <= "00000000";
--            LineBuffer1(1679) <= "00000000";
--            LineBuffer1(1680) <= "00000000";
--            LineBuffer1(1681) <= "00000000";
--            LineBuffer1(1682) <= "00000000";
--            LineBuffer1(1683) <= "00000000";
--            LineBuffer1(1684) <= "00000000";
--            LineBuffer1(1685) <= "00000000";
--            LineBuffer1(1686) <= "00000000";
--            LineBuffer1(1687) <= "00000000";
--            LineBuffer1(1688) <= "00000000";
--            LineBuffer1(1689) <= "00000000";    
--            LineBuffer1(1690) <= "00000000";
--            LineBuffer1(1691) <= "00000000";
--            LineBuffer1(1692) <= "00000000";
--            LineBuffer1(1693) <= "00000000";
--            LineBuffer1(1694) <= "00000000";
--            LineBuffer1(1695) <= "00000000";
--            LineBuffer1(1696) <= "00000000";
--            LineBuffer1(1697) <= "00000000";
--            LineBuffer1(1698) <= "00000000";
--            LineBuffer1(1699) <= "00000000";    
--            LineBuffer1(1700) <= "00000000";
--            LineBuffer1(1701) <= "00000000";
--            LineBuffer1(1702) <= "00000000";
--            LineBuffer1(1703) <= "00000000";
--            LineBuffer1(1704) <= "00000000";
--            LineBuffer1(1705) <= "00000000";
--            LineBuffer1(1706) <= "00000000";
--            LineBuffer1(1707) <= "00000000";
--            LineBuffer1(1708) <= "00000000";
--            LineBuffer1(1709) <= "00000000";    
--            LineBuffer1(1710) <= "00000000";
--            LineBuffer1(1711) <= "00000000";
--            LineBuffer1(1712) <= "00000000";
--            LineBuffer1(1713) <= "00000000";
--            LineBuffer1(1714) <= "00000000";
--            LineBuffer1(1715) <= "00000000";
--            LineBuffer1(1716) <= "00000000";
--            LineBuffer1(1717) <= "00000000";
--            LineBuffer1(1718) <= "00000000";
--            LineBuffer1(1719) <= "00000000";    
--            LineBuffer1(1720) <= "00000000";
--            LineBuffer1(1721) <= "00000000";
--            LineBuffer1(1722) <= "00000000";
--            LineBuffer1(1723) <= "00000000";
--            LineBuffer1(1724) <= "00000000";
--            LineBuffer1(1725) <= "00000000";
--            LineBuffer1(1726) <= "00000000";
--            LineBuffer1(1727) <= "00000000";
--            LineBuffer1(1728) <= "00000000";
--            LineBuffer1(1729) <= "00000000";    
--            LineBuffer1(1730) <= "00000000";
--            LineBuffer1(1731) <= "00000000";
--            LineBuffer1(1732) <= "00000000";
--            LineBuffer1(1733) <= "00000000";
--            LineBuffer1(1734) <= "00000000";
--            LineBuffer1(1735) <= "00000000";
--            LineBuffer1(1736) <= "00000000";
--            LineBuffer1(1737) <= "00000000";
--            LineBuffer1(1738) <= "00000000";
--            LineBuffer1(1739) <= "00000000";    
--            LineBuffer1(1740) <= "00000000";
--            LineBuffer1(1741) <= "00000000";
--            LineBuffer1(1742) <= "00000000";
--            LineBuffer1(1743) <= "00000000";
--            LineBuffer1(1744) <= "00000000";
--            LineBuffer1(1745) <= "00000000";
--            LineBuffer1(1746) <= "00000000";
--            LineBuffer1(1747) <= "00000000";
--            LineBuffer1(1748) <= "00000000";
--            LineBuffer1(1749) <= "00000000";    
--            LineBuffer1(1750) <= "00000000";
--            LineBuffer1(1751) <= "00000000";
--            LineBuffer1(1752) <= "00000000";
--            LineBuffer1(1753) <= "00000000";
--            LineBuffer1(1754) <= "00000000";
--            LineBuffer1(1755) <= "00000000";
--            LineBuffer1(1756) <= "00000000";
--            LineBuffer1(1757) <= "00000000";
--            LineBuffer1(1758) <= "00000000";
--            LineBuffer1(1759) <= "00000000";    
--            LineBuffer1(1760) <= "00000000";
--            LineBuffer1(1761) <= "00000000";
--            LineBuffer1(1762) <= "00000000";
--            LineBuffer1(1763) <= "00000000";
--            LineBuffer1(1764) <= "00000000";
--            LineBuffer1(1765) <= "00000000";
--            LineBuffer1(1766) <= "00000000";
--            LineBuffer1(1767) <= "00000000";
--            LineBuffer1(1768) <= "00000000";
--            LineBuffer1(1769) <= "00000000";    
--            LineBuffer1(1770) <= "00000000";
--            LineBuffer1(1771) <= "00000000";
--            LineBuffer1(1772) <= "00000000";
--            LineBuffer1(1773) <= "00000000";
--            LineBuffer1(1774) <= "00000000";
--            LineBuffer1(1775) <= "00000000";
--            LineBuffer1(1776) <= "00000000";
--            LineBuffer1(1777) <= "00000000";
--            LineBuffer1(1778) <= "00000000";
--            LineBuffer1(1779) <= "00000000";
--            LineBuffer1(1780) <= "00000000";
--            LineBuffer1(1781) <= "00000000";
--            LineBuffer1(1782) <= "00000000";
--            LineBuffer1(1783) <= "00000000";
--            LineBuffer1(1784) <= "00000000";
--            LineBuffer1(1785) <= "00000000";
--            LineBuffer1(1786) <= "00000000";
--            LineBuffer1(1787) <= "00000000";
--            LineBuffer1(1788) <= "00000000";
--            LineBuffer1(1789) <= "00000000";    
--            LineBuffer1(1790) <= "00000000";
--            LineBuffer1(1791) <= "00000000";
--            LineBuffer1(1792) <= "00000000";
--            LineBuffer1(1793) <= "00000000";
--            LineBuffer1(1794) <= "00000000";
--            LineBuffer1(1795) <= "00000000";
--            LineBuffer1(1796) <= "00000000";
--            LineBuffer1(1797) <= "00000000";
--            LineBuffer1(1798) <= "00000000";
--            LineBuffer1(1799) <= "00000000";    
--            LineBuffer1(1800) <= "00000000";
--            LineBuffer1(1801) <= "00000000";
--            LineBuffer1(1802) <= "00000000";
--            LineBuffer1(1803) <= "00000000";
--            LineBuffer1(1804) <= "00000000";
--            LineBuffer1(1805) <= "00000000";
--            LineBuffer1(1806) <= "00000000";
--            LineBuffer1(1807) <= "00000000";
--            LineBuffer1(1808) <= "00000000";
--            LineBuffer1(1809) <= "00000000";    
--            LineBuffer1(1810) <= "00000000";
--            LineBuffer1(1811) <= "00000000";
--            LineBuffer1(1812) <= "00000000";
--            LineBuffer1(1813) <= "00000000";
--            LineBuffer1(1814) <= "00000000";
--            LineBuffer1(1815) <= "00000000";
--            LineBuffer1(1816) <= "00000000";
--            LineBuffer1(1817) <= "00000000";
--            LineBuffer1(1818) <= "00000000";
--            LineBuffer1(1819) <= "00000000";    
--            LineBuffer1(1820) <= "00000000";
--            LineBuffer1(1821) <= "00000000";
--            LineBuffer1(1822) <= "00000000";
--            LineBuffer1(1823) <= "00000000";
--            LineBuffer1(1824) <= "00000000";
--            LineBuffer1(1825) <= "00000000";
--            LineBuffer1(1826) <= "00000000";
--            LineBuffer1(1827) <= "00000000";
--            LineBuffer1(1828) <= "00000000";
--            LineBuffer1(1829) <= "00000000";    
--            LineBuffer1(1830) <= "00000000";
--            LineBuffer1(1831) <= "00000000";
--            LineBuffer1(1832) <= "00000000";
--            LineBuffer1(1833) <= "00000000";
--            LineBuffer1(1834) <= "00000000";
--            LineBuffer1(1835) <= "00000000";
--            LineBuffer1(1836) <= "00000000";
--            LineBuffer1(1837) <= "00000000";
--            LineBuffer1(1838) <= "00000000";
--            LineBuffer1(1839) <= "00000000";    
--            LineBuffer1(1840) <= "00000000";
--            LineBuffer1(1841) <= "00000000";
--            LineBuffer1(1842) <= "00000000";
--            LineBuffer1(1843) <= "00000000";
--            LineBuffer1(1844) <= "00000000";
--            LineBuffer1(1845) <= "00000000";
--            LineBuffer1(1846) <= "00000000";
--            LineBuffer1(1847) <= "00000000";
--            LineBuffer1(1848) <= "00000000";
--            LineBuffer1(1849) <= "00000000";    
--            LineBuffer1(1850) <= "00000000";
--            LineBuffer1(1851) <= "00000000";
--            LineBuffer1(1852) <= "00000000";
--            LineBuffer1(1853) <= "00000000";
--            LineBuffer1(1854) <= "00000000";
--            LineBuffer1(1855) <= "00000000";
--            LineBuffer1(1856) <= "00000000";
--            LineBuffer1(1857) <= "00000000";
--            LineBuffer1(1858) <= "00000000";
--            LineBuffer1(1859) <= "00000000";    
--            LineBuffer1(1860) <= "00000000";
--            LineBuffer1(1861) <= "00000000";
--            LineBuffer1(1862) <= "00000000";
--            LineBuffer1(1863) <= "00000000";
--            LineBuffer1(1864) <= "00000000";
--            LineBuffer1(1865) <= "00000000";
--            LineBuffer1(1866) <= "00000000";
--            LineBuffer1(1867) <= "00000000";
--            LineBuffer1(1868) <= "00000000";
--            LineBuffer1(1869) <= "00000000";    
--            LineBuffer1(1870) <= "00000000";
--            LineBuffer1(1871) <= "00000000";
--            LineBuffer1(1872) <= "00000000";
--            LineBuffer1(1873) <= "00000000";
--            LineBuffer1(1874) <= "00000000";
--            LineBuffer1(1875) <= "00000000";
--            LineBuffer1(1876) <= "00000000";
--            LineBuffer1(1877) <= "00000000";
--            LineBuffer1(1878) <= "00000000";
--            LineBuffer1(1879) <= "00000000";
--            LineBuffer1(1880) <= "00000000";
--            LineBuffer1(1881) <= "00000000";
--            LineBuffer1(1882) <= "00000000";
--            LineBuffer1(1883) <= "00000000";
--            LineBuffer1(1884) <= "00000000";
--            LineBuffer1(1885) <= "00000000";
--            LineBuffer1(1886) <= "00000000";
--            LineBuffer1(1887) <= "00000000";
--            LineBuffer1(1888) <= "00000000";
--            LineBuffer1(1889) <= "00000000";    
--            LineBuffer1(1890) <= "00000000";
--            LineBuffer1(1891) <= "00000000";
--            LineBuffer1(1892) <= "00000000";
--            LineBuffer1(1893) <= "00000000";
--            LineBuffer1(1894) <= "00000000";
--            LineBuffer1(1895) <= "00000000";
--            LineBuffer1(1896) <= "00000000";
--            LineBuffer1(1897) <= "00000000";
--            LineBuffer1(1898) <= "00000000";
--            LineBuffer1(1899) <= "00000000";    
--            LineBuffer1(1900) <= "00000000";
--            LineBuffer1(1901) <= "00000000";
--            LineBuffer1(1902) <= "00000000";
--            LineBuffer1(1903) <= "00000000";
--            LineBuffer1(1904) <= "00000000";
--            LineBuffer1(1905) <= "00000000";
--            LineBuffer1(1906) <= "00000000";
--            LineBuffer1(1907) <= "00000000";
--            LineBuffer1(1908) <= "00000000";
--            LineBuffer1(1909) <= "00000000";    
--            LineBuffer1(1910) <= "00000000";
--            LineBuffer1(1911) <= "00000000";
--            LineBuffer1(1912) <= "00000000";
--            LineBuffer1(1913) <= "00000000";
--            LineBuffer1(1914) <= "00000000";
--            LineBuffer1(1915) <= "00000000";
--            LineBuffer1(1916) <= "00000000";
--            LineBuffer1(1917) <= "00000000";
--            LineBuffer1(1918) <= "00000000";
--            LineBuffer1(1919) <= "00000000";			
			
			
			
			
			
					
			LineBuffer2(0) <= "00000000";
			LineBuffer2(1) <= "00000000";
			LineBuffer2(2) <= "00000000";
			LineBuffer2(3) <= "00000000";
			LineBuffer2(4) <= "00000000";
			LineBuffer2(5) <= "00000000";
			LineBuffer2(6) <= "00000000";
			LineBuffer2(7) <= "00000000";
			LineBuffer2(8) <= "00000000";
			LineBuffer2(9) <= "00000000";	
			LineBuffer2(10) <= "00000000";
			LineBuffer2(11) <= "00000000";
			LineBuffer2(12) <= "00000000";
			LineBuffer2(13) <= "00000000";
			LineBuffer2(14) <= "00000000";
			LineBuffer2(15) <= "00000000";
			LineBuffer2(16) <= "00000000";
			LineBuffer2(17) <= "00000000";
			LineBuffer2(18) <= "00000000";
			LineBuffer2(19) <= "00000000";	
			LineBuffer2(20) <= "00000000";
			LineBuffer2(21) <= "00000000";
			LineBuffer2(22) <= "00000000";
			LineBuffer2(23) <= "00000000";
			LineBuffer2(24) <= "00000000";
			LineBuffer2(25) <= "00000000";
			LineBuffer2(26) <= "00000000";
			LineBuffer2(27) <= "00000000";
			LineBuffer2(28) <= "00000000";
			LineBuffer2(29) <= "00000000";	
			LineBuffer2(30) <= "00000000";
			LineBuffer2(31) <= "00000000";
			LineBuffer2(32) <= "00000000";
			LineBuffer2(33) <= "00000000";
			LineBuffer2(34) <= "00000000";
			LineBuffer2(35) <= "00000000";
			LineBuffer2(36) <= "00000000";
			LineBuffer2(37) <= "00000000";
			LineBuffer2(38) <= "00000000";
			LineBuffer2(39) <= "00000000";	
			LineBuffer2(40) <= "00000000";
			LineBuffer2(41) <= "00000000";
			LineBuffer2(42) <= "00000000";
			LineBuffer2(43) <= "00000000";
			LineBuffer2(44) <= "00000000";
			LineBuffer2(45) <= "00000000";
			LineBuffer2(46) <= "00000000";
			LineBuffer2(47) <= "00000000";
			LineBuffer2(48) <= "00000000";
			LineBuffer2(49) <= "00000000";	
			LineBuffer2(50) <= "00000000";
			LineBuffer2(51) <= "00000000";
			LineBuffer2(52) <= "00000000";
			LineBuffer2(53) <= "00000000";
			LineBuffer2(54) <= "00000000";
			LineBuffer2(55) <= "00000000";
			LineBuffer2(56) <= "00000000";
			LineBuffer2(57) <= "00000000";
			LineBuffer2(58) <= "00000000";
			LineBuffer2(59) <= "00000000";	
			LineBuffer2(60) <= "00000000";
			LineBuffer2(61) <= "00000000";
			LineBuffer2(62) <= "00000000";
			LineBuffer2(63) <= "00000000";
			LineBuffer2(64) <= "00000000";
			LineBuffer2(65) <= "00000000";
			LineBuffer2(66) <= "00000000";
			LineBuffer2(67) <= "00000000";
			LineBuffer2(68) <= "00000000";
			LineBuffer2(69) <= "00000000";	
			LineBuffer2(70) <= "00000000";
			LineBuffer2(71) <= "00000000";
			LineBuffer2(72) <= "00000000";
			LineBuffer2(73) <= "00000000";
			LineBuffer2(74) <= "00000000";
			LineBuffer2(75) <= "00000000";
			LineBuffer2(76) <= "00000000";
			LineBuffer2(77) <= "00000000";
			LineBuffer2(78) <= "00000000";
			LineBuffer2(79) <= "00000000";	
			LineBuffer2(80) <= "00000000";
			LineBuffer2(81) <= "00000000";
			LineBuffer2(82) <= "00000000";
			LineBuffer2(83) <= "00000000";
			LineBuffer2(84) <= "00000000";
			LineBuffer2(85) <= "00000000";
			LineBuffer2(86) <= "00000000";
			LineBuffer2(87) <= "00000000";
			LineBuffer2(88) <= "00000000";
			LineBuffer2(89) <= "00000000";	
			LineBuffer2(90) <= "00000000";
			LineBuffer2(91) <= "00000000";
			LineBuffer2(92) <= "00000000";
			LineBuffer2(93) <= "00000000";
			LineBuffer2(94) <= "00000000";
			LineBuffer2(95) <= "00000000";
			LineBuffer2(96) <= "00000000";
			LineBuffer2(97) <= "00000000";
			LineBuffer2(98) <= "00000000";
			LineBuffer2(99) <= "00000000";	
			LineBuffer2(100) <= "00000000";
			LineBuffer2(101) <= "00000000";
			LineBuffer2(102) <= "00000000";
			LineBuffer2(103) <= "00000000";
			LineBuffer2(104) <= "00000000";
			LineBuffer2(105) <= "00000000";
			LineBuffer2(106) <= "00000000";
			LineBuffer2(107) <= "00000000";
			LineBuffer2(108) <= "00000000";
			LineBuffer2(109) <= "00000000";	
			LineBuffer2(110) <= "00000000";
			LineBuffer2(111) <= "00000000";
			LineBuffer2(112) <= "00000000";
			LineBuffer2(113) <= "00000000";
			LineBuffer2(114) <= "00000000";
			LineBuffer2(115) <= "00000000";
			LineBuffer2(116) <= "00000000";
			LineBuffer2(117) <= "00000000";
			LineBuffer2(118) <= "00000000";
			LineBuffer2(119) <= "00000000";	
			LineBuffer2(120) <= "00000000";
			LineBuffer2(121) <= "00000000";
			LineBuffer2(122) <= "00000000";
			LineBuffer2(123) <= "00000000";
			LineBuffer2(124) <= "00000000";
			LineBuffer2(125) <= "00000000";
			LineBuffer2(126) <= "00000000";
			LineBuffer2(127) <= "00000000";
			LineBuffer2(128) <= "00000000";
			LineBuffer2(129) <= "00000000";	
			LineBuffer2(130) <= "00000000";
			LineBuffer2(131) <= "00000000";
			LineBuffer2(132) <= "00000000";
			LineBuffer2(133) <= "00000000";
			LineBuffer2(134) <= "00000000";
			LineBuffer2(135) <= "00000000";
			LineBuffer2(136) <= "00000000";
			LineBuffer2(137) <= "00000000";
			LineBuffer2(138) <= "00000000";
			LineBuffer2(139) <= "00000000";	
			LineBuffer2(140) <= "00000000";
			LineBuffer2(141) <= "00000000";
			LineBuffer2(142) <= "00000000";
			LineBuffer2(143) <= "00000000";
			LineBuffer2(144) <= "00000000";
			LineBuffer2(145) <= "00000000";
			LineBuffer2(146) <= "00000000";
			LineBuffer2(147) <= "00000000";
			LineBuffer2(148) <= "00000000";
			LineBuffer2(149) <= "00000000";	
			LineBuffer2(150) <= "00000000";
			LineBuffer2(151) <= "00000000";
			LineBuffer2(152) <= "00000000";
			LineBuffer2(153) <= "00000000";
			LineBuffer2(154) <= "00000000";
			LineBuffer2(155) <= "00000000";
			LineBuffer2(156) <= "00000000";
			LineBuffer2(157) <= "00000000";
			LineBuffer2(158) <= "00000000";
			LineBuffer2(159) <= "00000000";	
			LineBuffer2(160) <= "00000000";
			LineBuffer2(161) <= "00000000";
			LineBuffer2(162) <= "00000000";
			LineBuffer2(163) <= "00000000";
			LineBuffer2(164) <= "00000000";
			LineBuffer2(165) <= "00000000";
			LineBuffer2(166) <= "00000000";
			LineBuffer2(167) <= "00000000";
			LineBuffer2(168) <= "00000000";
			LineBuffer2(169) <= "00000000";	
			LineBuffer2(170) <= "00000000";
			LineBuffer2(171) <= "00000000";
			LineBuffer2(172) <= "00000000";
			LineBuffer2(173) <= "00000000";
			LineBuffer2(174) <= "00000000";
			LineBuffer2(175) <= "00000000";
			LineBuffer2(176) <= "00000000";
			LineBuffer2(177) <= "00000000";
			LineBuffer2(178) <= "00000000";
			LineBuffer2(179) <= "00000000";	
			LineBuffer2(180) <= "00000000";
			LineBuffer2(181) <= "00000000";
			LineBuffer2(182) <= "00000000";
			LineBuffer2(183) <= "00000000";
			LineBuffer2(184) <= "00000000";
			LineBuffer2(185) <= "00000000";
			LineBuffer2(186) <= "00000000";
			LineBuffer2(187) <= "00000000";
			LineBuffer2(188) <= "00000000";
			LineBuffer2(189) <= "00000000";	
			LineBuffer2(190) <= "00000000";
			LineBuffer2(191) <= "00000000";
			LineBuffer2(192) <= "00000000";
			LineBuffer2(193) <= "00000000";
			LineBuffer2(194) <= "00000000";
			LineBuffer2(195) <= "00000000";
			LineBuffer2(196) <= "00000000";
			LineBuffer2(197) <= "00000000";
			LineBuffer2(198) <= "00000000";
			LineBuffer2(199) <= "00000000";
			LineBuffer2(200) <= "00000000";
			LineBuffer2(201) <= "00000000";
			LineBuffer2(202) <= "00000000";
			LineBuffer2(203) <= "00000000";
			LineBuffer2(204) <= "00000000";
			LineBuffer2(205) <= "00000000";
			LineBuffer2(206) <= "00000000";
			LineBuffer2(207) <= "00000000";
			LineBuffer2(208) <= "00000000";
			LineBuffer2(209) <= "00000000";	
			LineBuffer2(210) <= "00000000";
			LineBuffer2(211) <= "00000000";
			LineBuffer2(212) <= "00000000";
			LineBuffer2(213) <= "00000000";
			LineBuffer2(214) <= "00000000";
			LineBuffer2(215) <= "00000000";
			LineBuffer2(216) <= "00000000";
			LineBuffer2(217) <= "00000000";
			LineBuffer2(218) <= "00000000";
			LineBuffer2(219) <= "00000000";	
			LineBuffer2(220) <= "00000000";
			LineBuffer2(221) <= "00000000";
			LineBuffer2(222) <= "00000000";
			LineBuffer2(223) <= "00000000";
			LineBuffer2(224) <= "00000000";
			LineBuffer2(225) <= "00000000";
			LineBuffer2(226) <= "00000000";
			LineBuffer2(227) <= "00000000";
			LineBuffer2(228) <= "00000000";
			LineBuffer2(229) <= "00000000";	
			LineBuffer2(230) <= "00000000";
			LineBuffer2(231) <= "00000000";
			LineBuffer2(232) <= "00000000";
			LineBuffer2(233) <= "00000000";
			LineBuffer2(234) <= "00000000";
			LineBuffer2(235) <= "00000000";
			LineBuffer2(236) <= "00000000";
			LineBuffer2(237) <= "00000000";
			LineBuffer2(238) <= "00000000";
			LineBuffer2(239) <= "00000000";	
			LineBuffer2(240) <= "00000000";
			LineBuffer2(241) <= "00000000";
			LineBuffer2(242) <= "00000000";
			LineBuffer2(243) <= "00000000";
			LineBuffer2(244) <= "00000000";
			LineBuffer2(245) <= "00000000";
			LineBuffer2(246) <= "00000000";
			LineBuffer2(247) <= "00000000";
			LineBuffer2(248) <= "00000000";
			LineBuffer2(249) <= "00000000";	
			LineBuffer2(250) <= "00000000";
			LineBuffer2(251) <= "00000000";
			LineBuffer2(252) <= "00000000";
			LineBuffer2(253) <= "00000000";
			LineBuffer2(254) <= "00000000";
			LineBuffer2(255) <= "00000000";
			LineBuffer2(256) <= "00000000";
			LineBuffer2(257) <= "00000000";
			LineBuffer2(258) <= "00000000";
			LineBuffer2(259) <= "00000000";	
			LineBuffer2(260) <= "00000000";
			LineBuffer2(261) <= "00000000";
			LineBuffer2(262) <= "00000000";
			LineBuffer2(263) <= "00000000";
			LineBuffer2(264) <= "00000000";
			LineBuffer2(265) <= "00000000";
			LineBuffer2(266) <= "00000000";
			LineBuffer2(267) <= "00000000";
			LineBuffer2(268) <= "00000000";
			LineBuffer2(269) <= "00000000";	
			LineBuffer2(270) <= "00000000";
			LineBuffer2(271) <= "00000000";
			LineBuffer2(272) <= "00000000";
			LineBuffer2(273) <= "00000000";
			LineBuffer2(274) <= "00000000";
			LineBuffer2(275) <= "00000000";
			LineBuffer2(276) <= "00000000";
			LineBuffer2(277) <= "00000000";
			LineBuffer2(278) <= "00000000";
			LineBuffer2(279) <= "00000000";	
			LineBuffer2(280) <= "00000000";
			LineBuffer2(281) <= "00000000";
			LineBuffer2(282) <= "00000000";
			LineBuffer2(283) <= "00000000";
			LineBuffer2(284) <= "00000000";
			LineBuffer2(285) <= "00000000";
			LineBuffer2(286) <= "00000000";
			LineBuffer2(287) <= "00000000";
			LineBuffer2(288) <= "00000000";
			LineBuffer2(289) <= "00000000";	
			LineBuffer2(290) <= "00000000";
			LineBuffer2(291) <= "00000000";
			LineBuffer2(292) <= "00000000";
			LineBuffer2(293) <= "00000000";
			LineBuffer2(294) <= "00000000";
			LineBuffer2(295) <= "00000000";
			LineBuffer2(296) <= "00000000";
			LineBuffer2(297) <= "00000000";
			LineBuffer2(298) <= "00000000";
			LineBuffer2(299) <= "00000000";
			LineBuffer2(300) <= "00000000";
			LineBuffer2(301) <= "00000000";
			LineBuffer2(302) <= "00000000";
			LineBuffer2(303) <= "00000000";
			LineBuffer2(304) <= "00000000";
			LineBuffer2(305) <= "00000000";
			LineBuffer2(306) <= "00000000";
			LineBuffer2(307) <= "00000000";
			LineBuffer2(308) <= "00000000";
			LineBuffer2(309) <= "00000000";	
			LineBuffer2(310) <= "00000000";
			LineBuffer2(311) <= "00000000";
			LineBuffer2(312) <= "00000000";
			LineBuffer2(313) <= "00000000";
			LineBuffer2(314) <= "00000000";
			LineBuffer2(315) <= "00000000";
			LineBuffer2(316) <= "00000000";
			LineBuffer2(317) <= "00000000";
			LineBuffer2(318) <= "00000000";
			LineBuffer2(319) <= "00000000";	
			LineBuffer2(320) <= "00000000";
			LineBuffer2(321) <= "00000000";
			LineBuffer2(322) <= "00000000";
			LineBuffer2(323) <= "00000000";
			LineBuffer2(324) <= "00000000";
			LineBuffer2(325) <= "00000000";
			LineBuffer2(326) <= "00000000";
			LineBuffer2(327) <= "00000000";
			LineBuffer2(328) <= "00000000";
			LineBuffer2(329) <= "00000000";	
			LineBuffer2(330) <= "00000000";
			LineBuffer2(331) <= "00000000";
			LineBuffer2(332) <= "00000000";
			LineBuffer2(333) <= "00000000";
			LineBuffer2(334) <= "00000000";
			LineBuffer2(335) <= "00000000";
			LineBuffer2(336) <= "00000000";
			LineBuffer2(337) <= "00000000";
			LineBuffer2(338) <= "00000000";
			LineBuffer2(339) <= "00000000";	
			LineBuffer2(340) <= "00000000";
			LineBuffer2(341) <= "00000000";
			LineBuffer2(342) <= "00000000";
			LineBuffer2(343) <= "00000000";
			LineBuffer2(344) <= "00000000";
			LineBuffer2(345) <= "00000000";
			LineBuffer2(346) <= "00000000";
			LineBuffer2(347) <= "00000000";
			LineBuffer2(348) <= "00000000";
			LineBuffer2(349) <= "00000000";	
			LineBuffer2(350) <= "00000000";
			LineBuffer2(351) <= "00000000";
			LineBuffer2(352) <= "00000000";
			LineBuffer2(353) <= "00000000";
			LineBuffer2(354) <= "00000000";
			LineBuffer2(355) <= "00000000";
			LineBuffer2(356) <= "00000000";
			LineBuffer2(357) <= "00000000";
			LineBuffer2(358) <= "00000000";
			LineBuffer2(359) <= "00000000";	
			LineBuffer2(360) <= "00000000";
			LineBuffer2(361) <= "00000000";
			LineBuffer2(362) <= "00000000";
			LineBuffer2(363) <= "00000000";
			LineBuffer2(364) <= "00000000";
			LineBuffer2(365) <= "00000000";
			LineBuffer2(366) <= "00000000";
			LineBuffer2(367) <= "00000000";
			LineBuffer2(368) <= "00000000";
			LineBuffer2(369) <= "00000000";	
			LineBuffer2(370) <= "00000000";
			LineBuffer2(371) <= "00000000";
			LineBuffer2(372) <= "00000000";
			LineBuffer2(373) <= "00000000";
			LineBuffer2(374) <= "00000000";
			LineBuffer2(375) <= "00000000";
			LineBuffer2(376) <= "00000000";
			LineBuffer2(377) <= "00000000";
			LineBuffer2(378) <= "00000000";
			LineBuffer2(379) <= "00000000";	
			LineBuffer2(380) <= "00000000";
			LineBuffer2(381) <= "00000000";
			LineBuffer2(382) <= "00000000";
			LineBuffer2(383) <= "00000000";
			LineBuffer2(384) <= "00000000";
			LineBuffer2(385) <= "00000000";
			LineBuffer2(386) <= "00000000";
			LineBuffer2(387) <= "00000000";
			LineBuffer2(388) <= "00000000";
			LineBuffer2(389) <= "00000000";	
			LineBuffer2(390) <= "00000000";
			LineBuffer2(391) <= "00000000";
			LineBuffer2(392) <= "00000000";
			LineBuffer2(393) <= "00000000";
			LineBuffer2(394) <= "00000000";
			LineBuffer2(395) <= "00000000";
			LineBuffer2(396) <= "00000000";
			LineBuffer2(397) <= "00000000";
			LineBuffer2(398) <= "00000000";
			LineBuffer2(399) <= "00000000";
			LineBuffer2(400) <= "00000000";
			LineBuffer2(401) <= "00000000";
			LineBuffer2(402) <= "00000000";
			LineBuffer2(403) <= "00000000";
			LineBuffer2(404) <= "00000000";
			LineBuffer2(405) <= "00000000";
			LineBuffer2(406) <= "00000000";
			LineBuffer2(407) <= "00000000";
			LineBuffer2(408) <= "00000000";
			LineBuffer2(409) <= "00000000";	
			LineBuffer2(410) <= "00000000";
			LineBuffer2(411) <= "00000000";
			LineBuffer2(412) <= "00000000";
			LineBuffer2(413) <= "00000000";
			LineBuffer2(414) <= "00000000";
			LineBuffer2(415) <= "00000000";
			LineBuffer2(416) <= "00000000";
			LineBuffer2(417) <= "00000000";
			LineBuffer2(418) <= "00000000";
			LineBuffer2(419) <= "00000000";	
			LineBuffer2(420) <= "00000000";
			LineBuffer2(421) <= "00000000";
			LineBuffer2(422) <= "00000000";
			LineBuffer2(423) <= "00000000";
			LineBuffer2(424) <= "00000000";
			LineBuffer2(425) <= "00000000";
			LineBuffer2(426) <= "00000000";
			LineBuffer2(427) <= "00000000";
			LineBuffer2(428) <= "00000000";
			LineBuffer2(429) <= "00000000";	
			LineBuffer2(430) <= "00000000";
			LineBuffer2(431) <= "00000000";
			LineBuffer2(432) <= "00000000";
			LineBuffer2(433) <= "00000000";
			LineBuffer2(434) <= "00000000";
			LineBuffer2(435) <= "00000000";
			LineBuffer2(436) <= "00000000";
			LineBuffer2(437) <= "00000000";
			LineBuffer2(438) <= "00000000";
			LineBuffer2(439) <= "00000000";	
			LineBuffer2(440) <= "00000000";
			LineBuffer2(441) <= "00000000";
			LineBuffer2(442) <= "00000000";
			LineBuffer2(443) <= "00000000";
			LineBuffer2(444) <= "00000000";
			LineBuffer2(445) <= "00000000";
			LineBuffer2(446) <= "00000000";
			LineBuffer2(447) <= "00000000";
			LineBuffer2(448) <= "00000000";
			LineBuffer2(449) <= "00000000";	
			LineBuffer2(450) <= "00000000";
			LineBuffer2(451) <= "00000000";
			LineBuffer2(452) <= "00000000";
			LineBuffer2(453) <= "00000000";
			LineBuffer2(454) <= "00000000";
			LineBuffer2(455) <= "00000000";
			LineBuffer2(456) <= "00000000";
			LineBuffer2(457) <= "00000000";
			LineBuffer2(458) <= "00000000";
			LineBuffer2(459) <= "00000000";	
			LineBuffer2(460) <= "00000000";
			LineBuffer2(461) <= "00000000";
			LineBuffer2(462) <= "00000000";
			LineBuffer2(463) <= "00000000";
			LineBuffer2(464) <= "00000000";
			LineBuffer2(465) <= "00000000";
			LineBuffer2(466) <= "00000000";
			LineBuffer2(467) <= "00000000";
			LineBuffer2(468) <= "00000000";
			LineBuffer2(469) <= "00000000";	
			LineBuffer2(470) <= "00000000";
			LineBuffer2(471) <= "00000000";
			LineBuffer2(472) <= "00000000";
			LineBuffer2(473) <= "00000000";
			LineBuffer2(474) <= "00000000";
			LineBuffer2(475) <= "00000000";
			LineBuffer2(476) <= "00000000";
			LineBuffer2(477) <= "00000000";
			LineBuffer2(478) <= "00000000";
			LineBuffer2(479) <= "00000000";	
			LineBuffer2(480) <= "00000000";
			LineBuffer2(481) <= "00000000";
			LineBuffer2(482) <= "00000000";
			LineBuffer2(483) <= "00000000";
			LineBuffer2(484) <= "00000000";
			LineBuffer2(485) <= "00000000";
			LineBuffer2(486) <= "00000000";
			LineBuffer2(487) <= "00000000";
			LineBuffer2(488) <= "00000000";
			LineBuffer2(489) <= "00000000";	
			LineBuffer2(490) <= "00000000";
			LineBuffer2(491) <= "00000000";
			LineBuffer2(492) <= "00000000";
			LineBuffer2(493) <= "00000000";
			LineBuffer2(494) <= "00000000";
			LineBuffer2(495) <= "00000000";
			LineBuffer2(496) <= "00000000";
			LineBuffer2(497) <= "00000000";
			LineBuffer2(498) <= "00000000";
			LineBuffer2(499) <= "00000000";
			LineBuffer2(500) <= "00000000";
			LineBuffer2(501) <= "00000000";
			LineBuffer2(502) <= "00000000";
			LineBuffer2(503) <= "00000000";
			LineBuffer2(504) <= "00000000";
			LineBuffer2(505) <= "00000000";
			LineBuffer2(506) <= "00000000";
			LineBuffer2(507) <= "00000000";
			LineBuffer2(508) <= "00000000";
			LineBuffer2(509) <= "00000000";	
			LineBuffer2(510) <= "00000000";
			LineBuffer2(511) <= "00000000";
			LineBuffer2(512) <= "00000000";
			LineBuffer2(513) <= "00000000";
			LineBuffer2(514) <= "00000000";
			LineBuffer2(515) <= "00000000";
			LineBuffer2(516) <= "00000000";
			LineBuffer2(517) <= "00000000";
			LineBuffer2(518) <= "00000000";
			LineBuffer2(519) <= "00000000";	
			LineBuffer2(520) <= "00000000";
			LineBuffer2(521) <= "00000000";
			LineBuffer2(522) <= "00000000";
			LineBuffer2(523) <= "00000000";
			LineBuffer2(524) <= "00000000";
			LineBuffer2(525) <= "00000000";
			LineBuffer2(526) <= "00000000";
			LineBuffer2(527) <= "00000000";
			LineBuffer2(528) <= "00000000";
			LineBuffer2(529) <= "00000000";	
			LineBuffer2(530) <= "00000000";
			LineBuffer2(531) <= "00000000";
			LineBuffer2(532) <= "00000000";
			LineBuffer2(533) <= "00000000";
			LineBuffer2(534) <= "00000000";
			LineBuffer2(535) <= "00000000";
			LineBuffer2(536) <= "00000000";
			LineBuffer2(537) <= "00000000";
			LineBuffer2(538) <= "00000000";
			LineBuffer2(539) <= "00000000";	
			LineBuffer2(540) <= "00000000";
			LineBuffer2(541) <= "00000000";
			LineBuffer2(542) <= "00000000";
			LineBuffer2(543) <= "00000000";
			LineBuffer2(544) <= "00000000";
			LineBuffer2(545) <= "00000000";
			LineBuffer2(546) <= "00000000";
			LineBuffer2(547) <= "00000000";
			LineBuffer2(548) <= "00000000";
			LineBuffer2(549) <= "00000000";	
			LineBuffer2(550) <= "00000000";
			LineBuffer2(551) <= "00000000";
			LineBuffer2(552) <= "00000000";
			LineBuffer2(553) <= "00000000";
			LineBuffer2(554) <= "00000000";
			LineBuffer2(555) <= "00000000";
			LineBuffer2(556) <= "00000000";
			LineBuffer2(557) <= "00000000";
			LineBuffer2(558) <= "00000000";
			LineBuffer2(559) <= "00000000";	
			LineBuffer2(560) <= "00000000";
			LineBuffer2(561) <= "00000000";
			LineBuffer2(562) <= "00000000";
			LineBuffer2(563) <= "00000000";
			LineBuffer2(564) <= "00000000";
			LineBuffer2(565) <= "00000000";
			LineBuffer2(566) <= "00000000";
			LineBuffer2(567) <= "00000000";
			LineBuffer2(568) <= "00000000";
			LineBuffer2(569) <= "00000000";	
			LineBuffer2(570) <= "00000000";
			LineBuffer2(571) <= "00000000";
			LineBuffer2(572) <= "00000000";
			LineBuffer2(573) <= "00000000";
			LineBuffer2(574) <= "00000000";
			LineBuffer2(575) <= "00000000";
			LineBuffer2(576) <= "00000000";
			LineBuffer2(577) <= "00000000";
			LineBuffer2(578) <= "00000000";
			LineBuffer2(579) <= "00000000";	
			LineBuffer2(580) <= "00000000";
			LineBuffer2(581) <= "00000000";
			LineBuffer2(582) <= "00000000";
			LineBuffer2(583) <= "00000000";
			LineBuffer2(584) <= "00000000";
			LineBuffer2(585) <= "00000000";
			LineBuffer2(586) <= "00000000";
			LineBuffer2(587) <= "00000000";
			LineBuffer2(588) <= "00000000";
			LineBuffer2(589) <= "00000000";	
			LineBuffer2(590) <= "00000000";
			LineBuffer2(591) <= "00000000";
			LineBuffer2(592) <= "00000000";
			LineBuffer2(593) <= "00000000";
			LineBuffer2(594) <= "00000000";
			LineBuffer2(595) <= "00000000";
			LineBuffer2(596) <= "00000000";
			LineBuffer2(597) <= "00000000";
			LineBuffer2(598) <= "00000000";
			LineBuffer2(599) <= "00000000";
			LineBuffer2(600) <= "00000000";
			LineBuffer2(601) <= "00000000";
			LineBuffer2(602) <= "00000000";
			LineBuffer2(603) <= "00000000";
			LineBuffer2(604) <= "00000000";
			LineBuffer2(605) <= "00000000";
			LineBuffer2(606) <= "00000000";
			LineBuffer2(607) <= "00000000";
			LineBuffer2(608) <= "00000000";
			LineBuffer2(609) <= "00000000";	
			LineBuffer2(610) <= "00000000";
			LineBuffer2(611) <= "00000000";
			LineBuffer2(612) <= "00000000";
			LineBuffer2(613) <= "00000000";
			LineBuffer2(614) <= "00000000";
			LineBuffer2(615) <= "00000000";
			LineBuffer2(616) <= "00000000";
			LineBuffer2(617) <= "00000000";
			LineBuffer2(618) <= "00000000";
			LineBuffer2(619) <= "00000000";	
			LineBuffer2(620) <= "00000000";
			LineBuffer2(621) <= "00000000";
			LineBuffer2(622) <= "00000000";
			LineBuffer2(623) <= "00000000";
			LineBuffer2(624) <= "00000000";
			LineBuffer2(625) <= "00000000";
			LineBuffer2(626) <= "00000000";
			LineBuffer2(627) <= "00000000";
			LineBuffer2(628) <= "00000000";
			LineBuffer2(629) <= "00000000";	
			LineBuffer2(630) <= "00000000";
			LineBuffer2(631) <= "00000000";
			LineBuffer2(632) <= "00000000";
			LineBuffer2(633) <= "00000000";
			LineBuffer2(634) <= "00000000";
			LineBuffer2(635) <= "00000000";
			LineBuffer2(636) <= "00000000";
			LineBuffer2(637) <= "00000000";
			LineBuffer2(638) <= "00000000";
			LineBuffer2(639) <= "00000000";
			LineBuffer2(640) <= "00000000";
            LineBuffer2(641) <= "00000000";
            LineBuffer2(642) <= "00000000";
            LineBuffer2(643) <= "00000000";
            LineBuffer2(644) <= "00000000";
            LineBuffer2(645) <= "00000000";
            LineBuffer2(646) <= "00000000";
            LineBuffer2(647) <= "00000000";
            LineBuffer2(648) <= "00000000";
            LineBuffer2(649) <= "00000000";    
            LineBuffer2(650) <= "00000000";
            LineBuffer2(651) <= "00000000";
            LineBuffer2(652) <= "00000000";
            LineBuffer2(653) <= "00000000";
            LineBuffer2(654) <= "00000000";
            LineBuffer2(655) <= "00000000";
            LineBuffer2(656) <= "00000000";
            LineBuffer2(657) <= "00000000";
            LineBuffer2(658) <= "00000000";
            LineBuffer2(659) <= "00000000";    
            LineBuffer2(660) <= "00000000";
            LineBuffer2(661) <= "00000000";
            LineBuffer2(662) <= "00000000";
            LineBuffer2(663) <= "00000000";
            LineBuffer2(664) <= "00000000";
            LineBuffer2(665) <= "00000000";
            LineBuffer2(666) <= "00000000";
            LineBuffer2(667) <= "00000000";
            LineBuffer2(668) <= "00000000";
            LineBuffer2(669) <= "00000000";    
            LineBuffer2(670) <= "00000000";
            LineBuffer2(671) <= "00000000";
            LineBuffer2(672) <= "00000000";
            LineBuffer2(673) <= "00000000";
            LineBuffer2(674) <= "00000000";
            LineBuffer2(675) <= "00000000";
            LineBuffer2(676) <= "00000000";
            LineBuffer2(677) <= "00000000";
            LineBuffer2(678) <= "00000000";
            LineBuffer2(679) <= "00000000";    
            LineBuffer2(680) <= "00000000";
            LineBuffer2(681) <= "00000000";
            LineBuffer2(682) <= "00000000";
            LineBuffer2(683) <= "00000000";
            LineBuffer2(684) <= "00000000";
            LineBuffer2(685) <= "00000000";
            LineBuffer2(686) <= "00000000";
            LineBuffer2(687) <= "00000000";
            LineBuffer2(688) <= "00000000";
            LineBuffer2(689) <= "00000000";    
            LineBuffer2(690) <= "00000000";
            LineBuffer2(691) <= "00000000";
            LineBuffer2(692) <= "00000000";
            LineBuffer2(693) <= "00000000";
            LineBuffer2(694) <= "00000000";
            LineBuffer2(695) <= "00000000";
            LineBuffer2(696) <= "00000000";
            LineBuffer2(697) <= "00000000";
            LineBuffer2(698) <= "00000000";
            LineBuffer2(699) <= "00000000";    
            LineBuffer2(700) <= "00000000";
            LineBuffer2(701) <= "00000000";
            LineBuffer2(702) <= "00000000";
            LineBuffer2(703) <= "00000000";
            LineBuffer2(704) <= "00000000";
            LineBuffer2(705) <= "00000000";
            LineBuffer2(706) <= "00000000";
            LineBuffer2(707) <= "00000000";
            LineBuffer2(708) <= "00000000";
            LineBuffer2(709) <= "00000000";    
            LineBuffer2(710) <= "00000000";
            LineBuffer2(711) <= "00000000";
            LineBuffer2(712) <= "00000000";
            LineBuffer2(713) <= "00000000";
            LineBuffer2(714) <= "00000000";
            LineBuffer2(715) <= "00000000";
            LineBuffer2(716) <= "00000000";
            LineBuffer2(717) <= "00000000";
            LineBuffer2(718) <= "00000000";
            LineBuffer2(719) <= "00000000";    
            LineBuffer2(720) <= "00000000";
            LineBuffer2(721) <= "00000000";
            LineBuffer2(722) <= "00000000";
            LineBuffer2(723) <= "00000000";
            LineBuffer2(724) <= "00000000";
            LineBuffer2(725) <= "00000000";
            LineBuffer2(726) <= "00000000";
            LineBuffer2(727) <= "00000000";
            LineBuffer2(728) <= "00000000";
            LineBuffer2(729) <= "00000000";    
            LineBuffer2(730) <= "00000000";
            LineBuffer2(731) <= "00000000";
            LineBuffer2(732) <= "00000000";
            LineBuffer2(733) <= "00000000";
            LineBuffer2(734) <= "00000000";
            LineBuffer2(735) <= "00000000";
            LineBuffer2(736) <= "00000000";
            LineBuffer2(737) <= "00000000";
            LineBuffer2(738) <= "00000000";
            LineBuffer2(739) <= "00000000";    
            LineBuffer2(740) <= "00000000";
            LineBuffer2(741) <= "00000000";
            LineBuffer2(742) <= "00000000";
            LineBuffer2(743) <= "00000000";
            LineBuffer2(744) <= "00000000";
            LineBuffer2(745) <= "00000000";
            LineBuffer2(746) <= "00000000";
            LineBuffer2(747) <= "00000000";
            LineBuffer2(748) <= "00000000";
            LineBuffer2(749) <= "00000000";    
            LineBuffer2(750) <= "00000000";
            LineBuffer2(751) <= "00000000";
            LineBuffer2(752) <= "00000000";
            LineBuffer2(753) <= "00000000";
            LineBuffer2(754) <= "00000000";
            LineBuffer2(755) <= "00000000";
            LineBuffer2(756) <= "00000000";
            LineBuffer2(757) <= "00000000";
            LineBuffer2(758) <= "00000000";
            LineBuffer2(759) <= "00000000";    
            LineBuffer2(760) <= "00000000";
            LineBuffer2(761) <= "00000000";
            LineBuffer2(762) <= "00000000";
            LineBuffer2(763) <= "00000000";
            LineBuffer2(764) <= "00000000";
            LineBuffer2(765) <= "00000000";
            LineBuffer2(766) <= "00000000";
            LineBuffer2(767) <= "00000000";
            LineBuffer2(768) <= "00000000";
            LineBuffer2(769) <= "00000000";    
            LineBuffer2(770) <= "00000000";
            LineBuffer2(771) <= "00000000";
            LineBuffer2(772) <= "00000000";
            LineBuffer2(773) <= "00000000";
            LineBuffer2(774) <= "00000000";
            LineBuffer2(775) <= "00000000";
            LineBuffer2(776) <= "00000000";
            LineBuffer2(777) <= "00000000";
            LineBuffer2(778) <= "00000000";
            LineBuffer2(779) <= "00000000";    
            LineBuffer2(780) <= "00000000";
            LineBuffer2(781) <= "00000000";
            LineBuffer2(782) <= "00000000";
            LineBuffer2(783) <= "00000000";
            LineBuffer2(784) <= "00000000";
            LineBuffer2(785) <= "00000000";
            LineBuffer2(786) <= "00000000";
            LineBuffer2(787) <= "00000000";
            LineBuffer2(788) <= "00000000";
            LineBuffer2(789) <= "00000000";    
            LineBuffer2(790) <= "00000000";
            LineBuffer2(791) <= "00000000";
            LineBuffer2(792) <= "00000000";
            LineBuffer2(793) <= "00000000";
            LineBuffer2(794) <= "00000000";
            LineBuffer2(795) <= "00000000";
            LineBuffer2(796) <= "00000000";
            LineBuffer2(797) <= "00000000";
            LineBuffer2(798) <= "00000000";
            LineBuffer2(799) <= "00000000";    
            LineBuffer2(800) <= "00000000";
            LineBuffer2(801) <= "00000000";
            LineBuffer2(802) <= "00000000";
            LineBuffer2(803) <= "00000000";
            LineBuffer2(804) <= "00000000";
            LineBuffer2(805) <= "00000000";
            LineBuffer2(806) <= "00000000";
            LineBuffer2(807) <= "00000000";
            LineBuffer2(808) <= "00000000";
            LineBuffer2(809) <= "00000000";    
            LineBuffer2(810) <= "00000000";
            LineBuffer2(811) <= "00000000";
            LineBuffer2(812) <= "00000000";
            LineBuffer2(813) <= "00000000";
            LineBuffer2(814) <= "00000000";
            LineBuffer2(815) <= "00000000";
            LineBuffer2(816) <= "00000000";
            LineBuffer2(817) <= "00000000";
            LineBuffer2(818) <= "00000000";
            LineBuffer2(819) <= "00000000";    
            LineBuffer2(820) <= "00000000";
            LineBuffer2(821) <= "00000000";
            LineBuffer2(822) <= "00000000";
            LineBuffer2(823) <= "00000000";
            LineBuffer2(824) <= "00000000";
            LineBuffer2(825) <= "00000000";
            LineBuffer2(826) <= "00000000";
            LineBuffer2(827) <= "00000000";
            LineBuffer2(828) <= "00000000";
            LineBuffer2(829) <= "00000000";    
            LineBuffer2(830) <= "00000000";
            LineBuffer2(831) <= "00000000";
            LineBuffer2(832) <= "00000000";
            LineBuffer2(833) <= "00000000";
            LineBuffer2(834) <= "00000000";
            LineBuffer2(835) <= "00000000";
            LineBuffer2(836) <= "00000000";
            LineBuffer2(837) <= "00000000";
            LineBuffer2(838) <= "00000000";
            LineBuffer2(839) <= "00000000";
            LineBuffer2(840) <= "00000000";
            LineBuffer2(841) <= "00000000";
            LineBuffer2(842) <= "00000000";
            LineBuffer2(843) <= "00000000";
            LineBuffer2(844) <= "00000000";
            LineBuffer2(845) <= "00000000";
            LineBuffer2(846) <= "00000000";
            LineBuffer2(847) <= "00000000";
            LineBuffer2(848) <= "00000000";
            LineBuffer2(849) <= "00000000";    
            LineBuffer2(850) <= "00000000";
            LineBuffer2(851) <= "00000000";
            LineBuffer2(852) <= "00000000";
            LineBuffer2(853) <= "00000000";
            LineBuffer2(854) <= "00000000";
            LineBuffer2(855) <= "00000000";
            LineBuffer2(856) <= "00000000";
            LineBuffer2(857) <= "00000000";
            LineBuffer2(858) <= "00000000";
            LineBuffer2(859) <= "00000000";    
            LineBuffer2(860) <= "00000000";
            LineBuffer2(861) <= "00000000";
            LineBuffer2(862) <= "00000000";
            LineBuffer2(863) <= "00000000";
            LineBuffer2(864) <= "00000000";
            LineBuffer2(865) <= "00000000";
            LineBuffer2(866) <= "00000000";
            LineBuffer2(867) <= "00000000";
            LineBuffer2(868) <= "00000000";
            LineBuffer2(869) <= "00000000";    
            LineBuffer2(870) <= "00000000";
            LineBuffer2(871) <= "00000000";
            LineBuffer2(872) <= "00000000";
            LineBuffer2(873) <= "00000000";
            LineBuffer2(874) <= "00000000";
            LineBuffer2(875) <= "00000000";
            LineBuffer2(876) <= "00000000";
            LineBuffer2(877) <= "00000000";
            LineBuffer2(878) <= "00000000";
            LineBuffer2(879) <= "00000000";    
            LineBuffer2(880) <= "00000000";
            LineBuffer2(881) <= "00000000";
            LineBuffer2(882) <= "00000000";
            LineBuffer2(883) <= "00000000";
            LineBuffer2(884) <= "00000000";
            LineBuffer2(885) <= "00000000";
            LineBuffer2(886) <= "00000000";
            LineBuffer2(887) <= "00000000";
            LineBuffer2(888) <= "00000000";
            LineBuffer2(889) <= "00000000";    
            LineBuffer2(890) <= "00000000";
            LineBuffer2(891) <= "00000000";
            LineBuffer2(892) <= "00000000";
            LineBuffer2(893) <= "00000000";
            LineBuffer2(894) <= "00000000";
            LineBuffer2(895) <= "00000000";
            LineBuffer2(896) <= "00000000";
            LineBuffer2(897) <= "00000000";
            LineBuffer2(898) <= "00000000";
            LineBuffer2(899) <= "00000000";    
            LineBuffer2(900) <= "00000000";
            LineBuffer2(901) <= "00000000";
            LineBuffer2(902) <= "00000000";
            LineBuffer2(903) <= "00000000";
            LineBuffer2(904) <= "00000000";
            LineBuffer2(905) <= "00000000";
            LineBuffer2(906) <= "00000000";
            LineBuffer2(907) <= "00000000";
            LineBuffer2(908) <= "00000000";
            LineBuffer2(909) <= "00000000";    
            LineBuffer2(910) <= "00000000";
            LineBuffer2(911) <= "00000000";
            LineBuffer2(912) <= "00000000";
            LineBuffer2(913) <= "00000000";
            LineBuffer2(914) <= "00000000";
            LineBuffer2(915) <= "00000000";
            LineBuffer2(916) <= "00000000";
            LineBuffer2(917) <= "00000000";
            LineBuffer2(918) <= "00000000";
            LineBuffer2(919) <= "00000000";    
            LineBuffer2(920) <= "00000000";
            LineBuffer2(921) <= "00000000";
            LineBuffer2(922) <= "00000000";
            LineBuffer2(923) <= "00000000";
            LineBuffer2(924) <= "00000000";
            LineBuffer2(925) <= "00000000";
            LineBuffer2(926) <= "00000000";
            LineBuffer2(927) <= "00000000";
            LineBuffer2(928) <= "00000000";
            LineBuffer2(929) <= "00000000";    
            LineBuffer2(930) <= "00000000";
            LineBuffer2(931) <= "00000000";
            LineBuffer2(932) <= "00000000";
            LineBuffer2(933) <= "00000000";
            LineBuffer2(934) <= "00000000";
            LineBuffer2(935) <= "00000000";
            LineBuffer2(936) <= "00000000";
            LineBuffer2(937) <= "00000000";
            LineBuffer2(938) <= "00000000";
            LineBuffer2(939) <= "00000000";
            LineBuffer2(940) <= "00000000";
            LineBuffer2(941) <= "00000000";
            LineBuffer2(942) <= "00000000";
            LineBuffer2(943) <= "00000000";
            LineBuffer2(944) <= "00000000";
            LineBuffer2(945) <= "00000000";
            LineBuffer2(946) <= "00000000";
            LineBuffer2(947) <= "00000000";
            LineBuffer2(948) <= "00000000";
            LineBuffer2(949) <= "00000000";    
            LineBuffer2(950) <= "00000000";
            LineBuffer2(951) <= "00000000";
            LineBuffer2(952) <= "00000000";
            LineBuffer2(953) <= "00000000";
            LineBuffer2(954) <= "00000000";
            LineBuffer2(955) <= "00000000";
            LineBuffer2(956) <= "00000000";
            LineBuffer2(957) <= "00000000";
            LineBuffer2(958) <= "00000000";
            LineBuffer2(959) <= "00000000";    
            LineBuffer2(960) <= "00000000";
            LineBuffer2(961) <= "00000000";
            LineBuffer2(962) <= "00000000";
            LineBuffer2(963) <= "00000000";
            LineBuffer2(964) <= "00000000";
            LineBuffer2(965) <= "00000000";
            LineBuffer2(966) <= "00000000";
            LineBuffer2(967) <= "00000000";
            LineBuffer2(968) <= "00000000";
            LineBuffer2(969) <= "00000000";    
            LineBuffer2(970) <= "00000000";
            LineBuffer2(971) <= "00000000";
            LineBuffer2(972) <= "00000000";
            LineBuffer2(973) <= "00000000";
            LineBuffer2(974) <= "00000000";
            LineBuffer2(975) <= "00000000";
            LineBuffer2(976) <= "00000000";
            LineBuffer2(977) <= "00000000";
            LineBuffer2(978) <= "00000000";
            LineBuffer2(979) <= "00000000";    
            LineBuffer2(980) <= "00000000";
            LineBuffer2(981) <= "00000000";
            LineBuffer2(982) <= "00000000";
            LineBuffer2(983) <= "00000000";
            LineBuffer2(984) <= "00000000";
            LineBuffer2(985) <= "00000000";
            LineBuffer2(986) <= "00000000";
            LineBuffer2(987) <= "00000000";
            LineBuffer2(988) <= "00000000";
            LineBuffer2(989) <= "00000000";    
            LineBuffer2(990) <= "00000000";
            LineBuffer2(991) <= "00000000";
            LineBuffer2(992) <= "00000000";
            LineBuffer2(993) <= "00000000";
            LineBuffer2(994) <= "00000000";
            LineBuffer2(995) <= "00000000";
            LineBuffer2(996) <= "00000000";
            LineBuffer2(997) <= "00000000";
            LineBuffer2(998) <= "00000000";
            LineBuffer2(999) <= "00000000";    
            LineBuffer2(1000) <= "00000000";
            LineBuffer2(1001) <= "00000000";
            LineBuffer2(1002) <= "00000000";
            LineBuffer2(1003) <= "00000000";
            LineBuffer2(1004) <= "00000000";
            LineBuffer2(1005) <= "00000000";
            LineBuffer2(1006) <= "00000000";
            LineBuffer2(1007) <= "00000000";
            LineBuffer2(1008) <= "00000000";
            LineBuffer2(1009) <= "00000000";    
            LineBuffer2(1010) <= "00000000";
            LineBuffer2(1011) <= "00000000";
            LineBuffer2(1012) <= "00000000";
            LineBuffer2(1013) <= "00000000";
            LineBuffer2(1014) <= "00000000";
            LineBuffer2(1015) <= "00000000";
            LineBuffer2(1016) <= "00000000";
            LineBuffer2(1017) <= "00000000";
            LineBuffer2(1018) <= "00000000";
            LineBuffer2(1019) <= "00000000";    
            LineBuffer2(1020) <= "00000000";
            LineBuffer2(1021) <= "00000000";
            LineBuffer2(1022) <= "00000000";
            LineBuffer2(1023) <= "00000000";
            LineBuffer2(1024) <= "00000000";
            LineBuffer2(1025) <= "00000000";
            LineBuffer2(1026) <= "00000000";
            LineBuffer2(1027) <= "00000000";
            LineBuffer2(1028) <= "00000000";
            LineBuffer2(1029) <= "00000000";    
            LineBuffer2(1030) <= "00000000";
            LineBuffer2(1031) <= "00000000";
            LineBuffer2(1032) <= "00000000";
            LineBuffer2(1033) <= "00000000";
            LineBuffer2(1034) <= "00000000";
            LineBuffer2(1035) <= "00000000";
            LineBuffer2(1036) <= "00000000";
            LineBuffer2(1037) <= "00000000";
            LineBuffer2(1038) <= "00000000";
            LineBuffer2(1039) <= "00000000";
            LineBuffer2(1040) <= "00000000";
            LineBuffer2(1041) <= "00000000";
            LineBuffer2(1042) <= "00000000";
            LineBuffer2(1043) <= "00000000";
            LineBuffer2(1044) <= "00000000";
            LineBuffer2(1045) <= "00000000";
            LineBuffer2(1046) <= "00000000";
            LineBuffer2(1047) <= "00000000";
            LineBuffer2(1048) <= "00000000";
            LineBuffer2(1049) <= "00000000";    
            LineBuffer2(1050) <= "00000000";
            LineBuffer2(1051) <= "00000000";
            LineBuffer2(1052) <= "00000000";
            LineBuffer2(1053) <= "00000000";
            LineBuffer2(1054) <= "00000000";
            LineBuffer2(1055) <= "00000000";
            LineBuffer2(1056) <= "00000000";
            LineBuffer2(1057) <= "00000000";
            LineBuffer2(1058) <= "00000000";
            LineBuffer2(1059) <= "00000000";    
            LineBuffer2(1060) <= "00000000";
            LineBuffer2(1061) <= "00000000";
            LineBuffer2(1062) <= "00000000";
            LineBuffer2(1063) <= "00000000";
            LineBuffer2(1064) <= "00000000";
            LineBuffer2(1065) <= "00000000";
            LineBuffer2(1066) <= "00000000";
            LineBuffer2(1067) <= "00000000";
            LineBuffer2(1068) <= "00000000";
            LineBuffer2(1069) <= "00000000";    
            LineBuffer2(1070) <= "00000000";
            LineBuffer2(1071) <= "00000000";
            LineBuffer2(1072) <= "00000000";
            LineBuffer2(1073) <= "00000000";
            LineBuffer2(1074) <= "00000000";
            LineBuffer2(1075) <= "00000000";
            LineBuffer2(1076) <= "00000000";
            LineBuffer2(1077) <= "00000000";
            LineBuffer2(1078) <= "00000000";
            LineBuffer2(1079) <= "00000000";    
            LineBuffer2(1080) <= "00000000";
            LineBuffer2(1081) <= "00000000";
            LineBuffer2(1082) <= "00000000";
            LineBuffer2(1083) <= "00000000";
            LineBuffer2(1084) <= "00000000";
            LineBuffer2(1085) <= "00000000";
            LineBuffer2(1086) <= "00000000";
            LineBuffer2(1087) <= "00000000";
            LineBuffer2(1088) <= "00000000";
            LineBuffer2(1089) <= "00000000";    
            LineBuffer2(1090) <= "00000000";
            LineBuffer2(1091) <= "00000000";
            LineBuffer2(1092) <= "00000000";
            LineBuffer2(1093) <= "00000000";
            LineBuffer2(1094) <= "00000000";
            LineBuffer2(1095) <= "00000000";
            LineBuffer2(1096) <= "00000000";
            LineBuffer2(1097) <= "00000000";
            LineBuffer2(1098) <= "00000000";
            LineBuffer2(1099) <= "00000000";    
            LineBuffer2(1100) <= "00000000";
            LineBuffer2(1101) <= "00000000";
            LineBuffer2(1102) <= "00000000";
            LineBuffer2(1103) <= "00000000";
            LineBuffer2(1104) <= "00000000";
            LineBuffer2(1105) <= "00000000";
            LineBuffer2(1106) <= "00000000";
            LineBuffer2(1107) <= "00000000";
            LineBuffer2(1108) <= "00000000";
            LineBuffer2(1109) <= "00000000";    
            LineBuffer2(1110) <= "00000000";
            LineBuffer2(1111) <= "00000000";
            LineBuffer2(1112) <= "00000000";
            LineBuffer2(1113) <= "00000000";
            LineBuffer2(1114) <= "00000000";
            LineBuffer2(1115) <= "00000000";
            LineBuffer2(1116) <= "00000000";
            LineBuffer2(1117) <= "00000000";
            LineBuffer2(1118) <= "00000000";
            LineBuffer2(1119) <= "00000000";    
            LineBuffer2(1120) <= "00000000";
            LineBuffer2(1121) <= "00000000";
            LineBuffer2(1122) <= "00000000";
            LineBuffer2(1123) <= "00000000";
            LineBuffer2(1124) <= "00000000";
            LineBuffer2(1125) <= "00000000";
            LineBuffer2(1126) <= "00000000";
            LineBuffer2(1127) <= "00000000";
            LineBuffer2(1128) <= "00000000";
            LineBuffer2(1129) <= "00000000";    
            LineBuffer2(1130) <= "00000000";
            LineBuffer2(1131) <= "00000000";
            LineBuffer2(1132) <= "00000000";
            LineBuffer2(1133) <= "00000000";
            LineBuffer2(1134) <= "00000000";
            LineBuffer2(1135) <= "00000000";
            LineBuffer2(1136) <= "00000000";
            LineBuffer2(1137) <= "00000000";
            LineBuffer2(1138) <= "00000000";
            LineBuffer2(1139) <= "00000000";
            LineBuffer2(1140) <= "00000000";
            LineBuffer2(1141) <= "00000000";
            LineBuffer2(1142) <= "00000000";
            LineBuffer2(1143) <= "00000000";
            LineBuffer2(1144) <= "00000000";
            LineBuffer2(1145) <= "00000000";
            LineBuffer2(1146) <= "00000000";
            LineBuffer2(1147) <= "00000000";
            LineBuffer2(1148) <= "00000000";
            LineBuffer2(1149) <= "00000000";    
            LineBuffer2(1150) <= "00000000";
            LineBuffer2(1151) <= "00000000";
            LineBuffer2(1152) <= "00000000";
            LineBuffer2(1153) <= "00000000";
            LineBuffer2(1154) <= "00000000";
            LineBuffer2(1155) <= "00000000";
            LineBuffer2(1156) <= "00000000";
            LineBuffer2(1157) <= "00000000";
            LineBuffer2(1158) <= "00000000";
            LineBuffer2(1159) <= "00000000";    
            LineBuffer2(1160) <= "00000000";
            LineBuffer2(1161) <= "00000000";
            LineBuffer2(1162) <= "00000000";
            LineBuffer2(1163) <= "00000000";
            LineBuffer2(1164) <= "00000000";
            LineBuffer2(1165) <= "00000000";
            LineBuffer2(1166) <= "00000000";
            LineBuffer2(1167) <= "00000000";
            LineBuffer2(1168) <= "00000000";
            LineBuffer2(1169) <= "00000000";    
            LineBuffer2(1170) <= "00000000";
            LineBuffer2(1171) <= "00000000";
            LineBuffer2(1172) <= "00000000";
            LineBuffer2(1173) <= "00000000";
            LineBuffer2(1174) <= "00000000";
            LineBuffer2(1175) <= "00000000";
            LineBuffer2(1176) <= "00000000";
            LineBuffer2(1177) <= "00000000";
            LineBuffer2(1178) <= "00000000";
            LineBuffer2(1179) <= "00000000";    
            LineBuffer2(1180) <= "00000000";
            LineBuffer2(1181) <= "00000000";
            LineBuffer2(1182) <= "00000000";
            LineBuffer2(1183) <= "00000000";
            LineBuffer2(1184) <= "00000000";
            LineBuffer2(1185) <= "00000000";
            LineBuffer2(1186) <= "00000000";
            LineBuffer2(1187) <= "00000000";
            LineBuffer2(1188) <= "00000000";
            LineBuffer2(1189) <= "00000000";    
            LineBuffer2(1190) <= "00000000";
            LineBuffer2(1191) <= "00000000";
            LineBuffer2(1192) <= "00000000";
            LineBuffer2(1193) <= "00000000";
            LineBuffer2(1194) <= "00000000";
            LineBuffer2(1195) <= "00000000";
            LineBuffer2(1196) <= "00000000";
            LineBuffer2(1197) <= "00000000";
            LineBuffer2(1198) <= "00000000";
            LineBuffer2(1199) <= "00000000";    
            LineBuffer2(1200) <= "00000000";
            LineBuffer2(1201) <= "00000000";
            LineBuffer2(1202) <= "00000000";
            LineBuffer2(1203) <= "00000000";
            LineBuffer2(1204) <= "00000000";
            LineBuffer2(1205) <= "00000000";
            LineBuffer2(1206) <= "00000000";
            LineBuffer2(1207) <= "00000000";
            LineBuffer2(1208) <= "00000000";
            LineBuffer2(1209) <= "00000000";    
            LineBuffer2(1210) <= "00000000";
            LineBuffer2(1211) <= "00000000";
            LineBuffer2(1212) <= "00000000";
            LineBuffer2(1213) <= "00000000";
            LineBuffer2(1214) <= "00000000";
            LineBuffer2(1215) <= "00000000";
            LineBuffer2(1216) <= "00000000";
            LineBuffer2(1217) <= "00000000";
            LineBuffer2(1218) <= "00000000";
            LineBuffer2(1219) <= "00000000";    
            LineBuffer2(1220) <= "00000000";
            LineBuffer2(1221) <= "00000000";
            LineBuffer2(1222) <= "00000000";
            LineBuffer2(1223) <= "00000000";
            LineBuffer2(1224) <= "00000000";
            LineBuffer2(1225) <= "00000000";
            LineBuffer2(1226) <= "00000000";
            LineBuffer2(1227) <= "00000000";
            LineBuffer2(1228) <= "00000000";
            LineBuffer2(1229) <= "00000000";    
            LineBuffer2(1230) <= "00000000";
            LineBuffer2(1231) <= "00000000";
            LineBuffer2(1232) <= "00000000";
            LineBuffer2(1233) <= "00000000";
            LineBuffer2(1234) <= "00000000";
            LineBuffer2(1235) <= "00000000";
            LineBuffer2(1236) <= "00000000";
            LineBuffer2(1237) <= "00000000";
            LineBuffer2(1238) <= "00000000";
            LineBuffer2(1239) <= "00000000";
            LineBuffer2(1240) <= "00000000";
            LineBuffer2(1241) <= "00000000";
            LineBuffer2(1242) <= "00000000";
            LineBuffer2(1243) <= "00000000";
            LineBuffer2(1244) <= "00000000";
            LineBuffer2(1245) <= "00000000";
            LineBuffer2(1246) <= "00000000";
            LineBuffer2(1247) <= "00000000";
            LineBuffer2(1248) <= "00000000";
            LineBuffer2(1249) <= "00000000";    
            LineBuffer2(1250) <= "00000000";
            LineBuffer2(1251) <= "00000000";
            LineBuffer2(1252) <= "00000000";
            LineBuffer2(1253) <= "00000000";
            LineBuffer2(1254) <= "00000000";
            LineBuffer2(1255) <= "00000000";
            LineBuffer2(1256) <= "00000000";
            LineBuffer2(1257) <= "00000000";
            LineBuffer2(1258) <= "00000000";
            LineBuffer2(1259) <= "00000000";    
            LineBuffer2(1260) <= "00000000";
            LineBuffer2(1261) <= "00000000";
            LineBuffer2(1262) <= "00000000";
            LineBuffer2(1263) <= "00000000";
            LineBuffer2(1264) <= "00000000";
            LineBuffer2(1265) <= "00000000";
            LineBuffer2(1266) <= "00000000";
            LineBuffer2(1267) <= "00000000";
            LineBuffer2(1268) <= "00000000";
            LineBuffer2(1269) <= "00000000";    
            LineBuffer2(1270) <= "00000000";
            LineBuffer2(1271) <= "00000000";
            LineBuffer2(1272) <= "00000000";
            LineBuffer2(1273) <= "00000000";
            LineBuffer2(1274) <= "00000000";
            LineBuffer2(1275) <= "00000000";
            LineBuffer2(1276) <= "00000000";
            LineBuffer2(1277) <= "00000000";
            LineBuffer2(1278) <= "00000000";
            LineBuffer2(1279) <= "00000000";
            
            
--            LineBuffer2(1280) <= "00000000";
--            LineBuffer2(1281) <= "00000000";
--            LineBuffer2(1282) <= "00000000";
--            LineBuffer2(1283) <= "00000000";
--            LineBuffer2(1284) <= "00000000";
--            LineBuffer2(1285) <= "00000000";
--            LineBuffer2(1286) <= "00000000";
--            LineBuffer2(1287) <= "00000000";
--            LineBuffer2(1288) <= "00000000";
--            LineBuffer2(1289) <= "00000000";    
--            LineBuffer2(1290) <= "00000000";
--            LineBuffer2(1291) <= "00000000";
--            LineBuffer2(1292) <= "00000000";
--            LineBuffer2(1293) <= "00000000";
--            LineBuffer2(1294) <= "00000000";
--            LineBuffer2(1295) <= "00000000";
--            LineBuffer2(1296) <= "00000000";
--            LineBuffer2(1297) <= "00000000";
--            LineBuffer2(1298) <= "00000000";
--            LineBuffer2(1299) <= "00000000";    
--            LineBuffer2(1300) <= "00000000";
--            LineBuffer2(1301) <= "00000000";
--            LineBuffer2(1302) <= "00000000";
--            LineBuffer2(1303) <= "00000000";
--            LineBuffer2(1304) <= "00000000";
--            LineBuffer2(1305) <= "00000000";
--            LineBuffer2(1306) <= "00000000";
--            LineBuffer2(1307) <= "00000000";
--            LineBuffer2(1308) <= "00000000";
--            LineBuffer2(1309) <= "00000000";    
--            LineBuffer2(1310) <= "00000000";
--            LineBuffer2(1311) <= "00000000";
--            LineBuffer2(1312) <= "00000000";
--            LineBuffer2(1313) <= "00000000";
--            LineBuffer2(1314) <= "00000000";
--            LineBuffer2(1315) <= "00000000";
--            LineBuffer2(1316) <= "00000000";
--            LineBuffer2(1317) <= "00000000";
--            LineBuffer2(1318) <= "00000000";
--            LineBuffer2(1319) <= "00000000";    
--            LineBuffer2(1320) <= "00000000";
--            LineBuffer2(1321) <= "00000000";
--            LineBuffer2(1322) <= "00000000";
--            LineBuffer2(1323) <= "00000000";
--            LineBuffer2(1324) <= "00000000";
--            LineBuffer2(1325) <= "00000000";
--            LineBuffer2(1326) <= "00000000";
--            LineBuffer2(1327) <= "00000000";
--            LineBuffer2(1328) <= "00000000";
--            LineBuffer2(1329) <= "00000000";    
--            LineBuffer2(1330) <= "00000000";
--            LineBuffer2(1331) <= "00000000";
--            LineBuffer2(1332) <= "00000000";
--            LineBuffer2(1333) <= "00000000";
--            LineBuffer2(1334) <= "00000000";
--            LineBuffer2(1335) <= "00000000";
--            LineBuffer2(1336) <= "00000000";
--            LineBuffer2(1337) <= "00000000";
--            LineBuffer2(1338) <= "00000000";
--            LineBuffer2(1339) <= "00000000";    
--            LineBuffer2(1340) <= "00000000";
--            LineBuffer2(1341) <= "00000000";
--            LineBuffer2(1342) <= "00000000";
--            LineBuffer2(1343) <= "00000000";
--            LineBuffer2(1344) <= "00000000";
--            LineBuffer2(1345) <= "00000000";
--            LineBuffer2(1346) <= "00000000";
--            LineBuffer2(1347) <= "00000000";
--            LineBuffer2(1348) <= "00000000";
--            LineBuffer2(1349) <= "00000000";    
--            LineBuffer2(1350) <= "00000000";
--            LineBuffer2(1351) <= "00000000";
--            LineBuffer2(1352) <= "00000000";
--            LineBuffer2(1353) <= "00000000";
--            LineBuffer2(1354) <= "00000000";
--            LineBuffer2(1355) <= "00000000";
--            LineBuffer2(1356) <= "00000000";
--            LineBuffer2(1357) <= "00000000";
--            LineBuffer2(1358) <= "00000000";
--            LineBuffer2(1359) <= "00000000";    
--            LineBuffer2(1360) <= "00000000";
--            LineBuffer2(1361) <= "00000000";
--            LineBuffer2(1362) <= "00000000";
--            LineBuffer2(1363) <= "00000000";
--            LineBuffer2(1364) <= "00000000";
--            LineBuffer2(1365) <= "00000000";
--            LineBuffer2(1366) <= "00000000";
--            LineBuffer2(1367) <= "00000000";
--            LineBuffer2(1368) <= "00000000";
--            LineBuffer2(1369) <= "00000000";    
--            LineBuffer2(1370) <= "00000000";
--            LineBuffer2(1371) <= "00000000";
--            LineBuffer2(1372) <= "00000000";
--            LineBuffer2(1373) <= "00000000";
--            LineBuffer2(1374) <= "00000000";
--            LineBuffer2(1375) <= "00000000";
--            LineBuffer2(1376) <= "00000000";
--            LineBuffer2(1377) <= "00000000";
--            LineBuffer2(1378) <= "00000000";
--            LineBuffer2(1379) <= "00000000";    
--            LineBuffer2(1380) <= "00000000";
--            LineBuffer2(1381) <= "00000000";
--            LineBuffer2(1382) <= "00000000";
--            LineBuffer2(1383) <= "00000000";
--            LineBuffer2(1384) <= "00000000";
--            LineBuffer2(1385) <= "00000000";
--            LineBuffer2(1386) <= "00000000";
--            LineBuffer2(1387) <= "00000000";
--            LineBuffer2(1388) <= "00000000";
--            LineBuffer2(1389) <= "00000000";    
--            LineBuffer2(1390) <= "00000000";
--            LineBuffer2(1391) <= "00000000";
--            LineBuffer2(1392) <= "00000000";
--            LineBuffer2(1393) <= "00000000";
--            LineBuffer2(1394) <= "00000000";
--            LineBuffer2(1395) <= "00000000";
--            LineBuffer2(1396) <= "00000000";
--            LineBuffer2(1397) <= "00000000";
--            LineBuffer2(1398) <= "00000000";
--            LineBuffer2(1399) <= "00000000";    
--            LineBuffer2(1400) <= "00000000";
--            LineBuffer2(1401) <= "00000000";
--            LineBuffer2(1402) <= "00000000";
--            LineBuffer2(1403) <= "00000000";
--            LineBuffer2(1404) <= "00000000";
--            LineBuffer2(1405) <= "00000000";
--            LineBuffer2(1406) <= "00000000";
--            LineBuffer2(1407) <= "00000000";
--            LineBuffer2(1408) <= "00000000";
--            LineBuffer2(1409) <= "00000000";    
--            LineBuffer2(1410) <= "00000000";
--            LineBuffer2(1411) <= "00000000";
--            LineBuffer2(1412) <= "00000000";
--            LineBuffer2(1413) <= "00000000";
--            LineBuffer2(1414) <= "00000000";
--            LineBuffer2(1415) <= "00000000";
--            LineBuffer2(1416) <= "00000000";
--            LineBuffer2(1417) <= "00000000";
--            LineBuffer2(1418) <= "00000000";
--            LineBuffer2(1419) <= "00000000";    
--            LineBuffer2(1420) <= "00000000";
--            LineBuffer2(1421) <= "00000000";
--            LineBuffer2(1422) <= "00000000";
--            LineBuffer2(1423) <= "00000000";
--            LineBuffer2(1424) <= "00000000";
--            LineBuffer2(1425) <= "00000000";
--            LineBuffer2(1426) <= "00000000";
--            LineBuffer2(1427) <= "00000000";
--            LineBuffer2(1428) <= "00000000";
--            LineBuffer2(1429) <= "00000000";    
--            LineBuffer2(1430) <= "00000000";
--            LineBuffer2(1431) <= "00000000";
--            LineBuffer2(1432) <= "00000000";
--            LineBuffer2(1433) <= "00000000";
--            LineBuffer2(1434) <= "00000000";
--            LineBuffer2(1435) <= "00000000";
--            LineBuffer2(1436) <= "00000000";
--            LineBuffer2(1437) <= "00000000";
--            LineBuffer2(1438) <= "00000000";
--            LineBuffer2(1439) <= "00000000";    
--            LineBuffer2(1440) <= "00000000";
--            LineBuffer2(1441) <= "00000000";
--            LineBuffer2(1442) <= "00000000";
--            LineBuffer2(1443) <= "00000000";
--            LineBuffer2(1444) <= "00000000";
--            LineBuffer2(1445) <= "00000000";
--            LineBuffer2(1446) <= "00000000";
--            LineBuffer2(1447) <= "00000000";
--            LineBuffer2(1448) <= "00000000";
--            LineBuffer2(1449) <= "00000000";    
--            LineBuffer2(1450) <= "00000000";
--            LineBuffer2(1451) <= "00000000";
--            LineBuffer2(1452) <= "00000000";
--            LineBuffer2(1453) <= "00000000";
--            LineBuffer2(1454) <= "00000000";
--            LineBuffer2(1455) <= "00000000";
--            LineBuffer2(1456) <= "00000000";
--            LineBuffer2(1457) <= "00000000";
--            LineBuffer2(1458) <= "00000000";
--            LineBuffer2(1459) <= "00000000";    
--            LineBuffer2(1460) <= "00000000";
--            LineBuffer2(1461) <= "00000000";
--            LineBuffer2(1462) <= "00000000";
--            LineBuffer2(1463) <= "00000000";
--            LineBuffer2(1464) <= "00000000";
--            LineBuffer2(1465) <= "00000000";
--            LineBuffer2(1466) <= "00000000";
--            LineBuffer2(1467) <= "00000000";
--            LineBuffer2(1468) <= "00000000";
--            LineBuffer2(1469) <= "00000000";    
--            LineBuffer2(1470) <= "00000000";
--            LineBuffer2(1471) <= "00000000";
--            LineBuffer2(1472) <= "00000000";
--            LineBuffer2(1473) <= "00000000";
--            LineBuffer2(1474) <= "00000000";
--            LineBuffer2(1475) <= "00000000";
--            LineBuffer2(1476) <= "00000000";
--            LineBuffer2(1477) <= "00000000";
--            LineBuffer2(1478) <= "00000000";
--            LineBuffer2(1479) <= "00000000";
--            LineBuffer2(1480) <= "00000000";
--            LineBuffer2(1481) <= "00000000";
--            LineBuffer2(1482) <= "00000000";
--            LineBuffer2(1483) <= "00000000";
--            LineBuffer2(1484) <= "00000000";
--            LineBuffer2(1485) <= "00000000";
--            LineBuffer2(1486) <= "00000000";
--            LineBuffer2(1487) <= "00000000";
--            LineBuffer2(1488) <= "00000000";
--            LineBuffer2(1489) <= "00000000";    
--            LineBuffer2(1490) <= "00000000";
--            LineBuffer2(1491) <= "00000000";
--            LineBuffer2(1492) <= "00000000";
--            LineBuffer2(1493) <= "00000000";
--            LineBuffer2(1494) <= "00000000";
--            LineBuffer2(1495) <= "00000000";
--            LineBuffer2(1496) <= "00000000";
--            LineBuffer2(1497) <= "00000000";
--            LineBuffer2(1498) <= "00000000";
--            LineBuffer2(1499) <= "00000000";    
--            LineBuffer2(1500) <= "00000000";
--            LineBuffer2(1501) <= "00000000";
--            LineBuffer2(1502) <= "00000000";
--            LineBuffer2(1503) <= "00000000";
--            LineBuffer2(1504) <= "00000000";
--            LineBuffer2(1505) <= "00000000";
--            LineBuffer2(1506) <= "00000000";
--            LineBuffer2(1507) <= "00000000";
--            LineBuffer2(1508) <= "00000000";
--            LineBuffer2(1509) <= "00000000";    
--            LineBuffer2(1510) <= "00000000";
--            LineBuffer2(1511) <= "00000000";
--            LineBuffer2(1512) <= "00000000";
--            LineBuffer2(1513) <= "00000000";
--            LineBuffer2(1514) <= "00000000";
--            LineBuffer2(1515) <= "00000000";
--            LineBuffer2(1516) <= "00000000";
--            LineBuffer2(1517) <= "00000000";
--            LineBuffer2(1518) <= "00000000";
--            LineBuffer2(1519) <= "00000000";    
--            LineBuffer2(1520) <= "00000000";
--            LineBuffer2(1521) <= "00000000";
--            LineBuffer2(1522) <= "00000000";
--            LineBuffer2(1523) <= "00000000";
--            LineBuffer2(1524) <= "00000000";
--            LineBuffer2(1525) <= "00000000";
--            LineBuffer2(1526) <= "00000000";
--            LineBuffer2(1527) <= "00000000";
--            LineBuffer2(1528) <= "00000000";
--            LineBuffer2(1529) <= "00000000";    
--            LineBuffer2(1530) <= "00000000";
--            LineBuffer2(1531) <= "00000000";
--            LineBuffer2(1532) <= "00000000";
--            LineBuffer2(1533) <= "00000000";
--            LineBuffer2(1534) <= "00000000";
--            LineBuffer2(1535) <= "00000000";
--            LineBuffer2(1536) <= "00000000";
--            LineBuffer2(1537) <= "00000000";
--            LineBuffer2(1538) <= "00000000";
--            LineBuffer2(1539) <= "00000000";    
--            LineBuffer2(1540) <= "00000000";
--            LineBuffer2(1541) <= "00000000";
--            LineBuffer2(1542) <= "00000000";
--            LineBuffer2(1543) <= "00000000";
--            LineBuffer2(1544) <= "00000000";
--            LineBuffer2(1545) <= "00000000";
--            LineBuffer2(1546) <= "00000000";
--            LineBuffer2(1547) <= "00000000";
--            LineBuffer2(1548) <= "00000000";
--            LineBuffer2(1549) <= "00000000";    
--            LineBuffer2(1550) <= "00000000";
--            LineBuffer2(1551) <= "00000000";
--            LineBuffer2(1552) <= "00000000";
--            LineBuffer2(1553) <= "00000000";
--            LineBuffer2(1554) <= "00000000";
--            LineBuffer2(1555) <= "00000000";
--            LineBuffer2(1556) <= "00000000";
--            LineBuffer2(1557) <= "00000000";
--            LineBuffer2(1558) <= "00000000";
--            LineBuffer2(1559) <= "00000000";    
--            LineBuffer2(1560) <= "00000000";
--            LineBuffer2(1561) <= "00000000";
--            LineBuffer2(1562) <= "00000000";
--            LineBuffer2(1563) <= "00000000";
--            LineBuffer2(1564) <= "00000000";
--            LineBuffer2(1565) <= "00000000";
--            LineBuffer2(1566) <= "00000000";
--            LineBuffer2(1567) <= "00000000";
--            LineBuffer2(1568) <= "00000000";
--            LineBuffer2(1569) <= "00000000";    
--            LineBuffer2(1570) <= "00000000";
--            LineBuffer2(1571) <= "00000000";
--            LineBuffer2(1572) <= "00000000";
--            LineBuffer2(1573) <= "00000000";
--            LineBuffer2(1574) <= "00000000";
--            LineBuffer2(1575) <= "00000000";
--            LineBuffer2(1576) <= "00000000";
--            LineBuffer2(1577) <= "00000000";
--            LineBuffer2(1578) <= "00000000";
--            LineBuffer2(1579) <= "00000000";
--            LineBuffer2(1580) <= "00000000";
--            LineBuffer2(1581) <= "00000000";
--            LineBuffer2(1582) <= "00000000";
--            LineBuffer2(1583) <= "00000000";
--            LineBuffer2(1584) <= "00000000";
--            LineBuffer2(1585) <= "00000000";
--            LineBuffer2(1586) <= "00000000";
--            LineBuffer2(1587) <= "00000000";
--            LineBuffer2(1588) <= "00000000";
--            LineBuffer2(1589) <= "00000000";    
--            LineBuffer2(1590) <= "00000000";
--            LineBuffer2(1591) <= "00000000";
--            LineBuffer2(1592) <= "00000000";
--            LineBuffer2(1593) <= "00000000";
--            LineBuffer2(1594) <= "00000000";
--            LineBuffer2(1595) <= "00000000";
--            LineBuffer2(1596) <= "00000000";
--            LineBuffer2(1597) <= "00000000";
--            LineBuffer2(1598) <= "00000000";
--            LineBuffer2(1599) <= "00000000";    
--            LineBuffer2(1600) <= "00000000";
--            LineBuffer2(1601) <= "00000000";
--            LineBuffer2(1602) <= "00000000";
--            LineBuffer2(1603) <= "00000000";
--            LineBuffer2(1604) <= "00000000";
--            LineBuffer2(1605) <= "00000000";
--            LineBuffer2(1606) <= "00000000";
--            LineBuffer2(1607) <= "00000000";
--            LineBuffer2(1608) <= "00000000";
--            LineBuffer2(1609) <= "00000000";    
--            LineBuffer2(1610) <= "00000000";
--            LineBuffer2(1611) <= "00000000";
--            LineBuffer2(1612) <= "00000000";
--            LineBuffer2(1613) <= "00000000";
--            LineBuffer2(1614) <= "00000000";
--            LineBuffer2(1615) <= "00000000";
--            LineBuffer2(1616) <= "00000000";
--            LineBuffer2(1617) <= "00000000";
--            LineBuffer2(1618) <= "00000000";
--            LineBuffer2(1619) <= "00000000";    
--            LineBuffer2(1620) <= "00000000";
--            LineBuffer2(1621) <= "00000000";
--            LineBuffer2(1622) <= "00000000";
--            LineBuffer2(1623) <= "00000000";
--            LineBuffer2(1624) <= "00000000";
--            LineBuffer2(1625) <= "00000000";
--            LineBuffer2(1626) <= "00000000";
--            LineBuffer2(1627) <= "00000000";
--            LineBuffer2(1628) <= "00000000";
--            LineBuffer2(1629) <= "00000000";    
--            LineBuffer2(1630) <= "00000000";
--            LineBuffer2(1631) <= "00000000";
--            LineBuffer2(1632) <= "00000000";
--            LineBuffer2(1633) <= "00000000";
--            LineBuffer2(1634) <= "00000000";
--            LineBuffer2(1635) <= "00000000";
--            LineBuffer2(1636) <= "00000000";
--            LineBuffer2(1637) <= "00000000";
--            LineBuffer2(1638) <= "00000000";
--            LineBuffer2(1639) <= "00000000";    
--            LineBuffer2(1640) <= "00000000";
--            LineBuffer2(1641) <= "00000000";
--            LineBuffer2(1642) <= "00000000";
--            LineBuffer2(1643) <= "00000000";
--            LineBuffer2(1644) <= "00000000";
--            LineBuffer2(1645) <= "00000000";
--            LineBuffer2(1646) <= "00000000";
--            LineBuffer2(1647) <= "00000000";
--            LineBuffer2(1648) <= "00000000";
--            LineBuffer2(1649) <= "00000000";    
--            LineBuffer2(1650) <= "00000000";
--            LineBuffer2(1651) <= "00000000";
--            LineBuffer2(1652) <= "00000000";
--            LineBuffer2(1653) <= "00000000";
--            LineBuffer2(1654) <= "00000000";
--            LineBuffer2(1655) <= "00000000";
--            LineBuffer2(1656) <= "00000000";
--            LineBuffer2(1657) <= "00000000";
--            LineBuffer2(1658) <= "00000000";
--            LineBuffer2(1659) <= "00000000";    
--            LineBuffer2(1660) <= "00000000";
--            LineBuffer2(1661) <= "00000000";
--            LineBuffer2(1662) <= "00000000";
--            LineBuffer2(1663) <= "00000000";
--            LineBuffer2(1664) <= "00000000";
--            LineBuffer2(1665) <= "00000000";
--            LineBuffer2(1666) <= "00000000";
--            LineBuffer2(1667) <= "00000000";
--            LineBuffer2(1668) <= "00000000";
--            LineBuffer2(1669) <= "00000000";    
--            LineBuffer2(1670) <= "00000000";
--            LineBuffer2(1671) <= "00000000";
--            LineBuffer2(1672) <= "00000000";
--            LineBuffer2(1673) <= "00000000";
--            LineBuffer2(1674) <= "00000000";
--            LineBuffer2(1675) <= "00000000";
--            LineBuffer2(1676) <= "00000000";
--            LineBuffer2(1677) <= "00000000";
--            LineBuffer2(1678) <= "00000000";
--            LineBuffer2(1679) <= "00000000";
--            LineBuffer2(1680) <= "00000000";
--            LineBuffer2(1681) <= "00000000";
--            LineBuffer2(1682) <= "00000000";
--            LineBuffer2(1683) <= "00000000";
--            LineBuffer2(1684) <= "00000000";
--            LineBuffer2(1685) <= "00000000";
--            LineBuffer2(1686) <= "00000000";
--            LineBuffer2(1687) <= "00000000";
--            LineBuffer2(1688) <= "00000000";
--            LineBuffer2(1689) <= "00000000";    
--            LineBuffer2(1690) <= "00000000";
--            LineBuffer2(1691) <= "00000000";
--            LineBuffer2(1692) <= "00000000";
--            LineBuffer2(1693) <= "00000000";
--            LineBuffer2(1694) <= "00000000";
--            LineBuffer2(1695) <= "00000000";
--            LineBuffer2(1696) <= "00000000";
--            LineBuffer2(1697) <= "00000000";
--            LineBuffer2(1698) <= "00000000";
--            LineBuffer2(1699) <= "00000000";    
--            LineBuffer2(1700) <= "00000000";
--            LineBuffer2(1701) <= "00000000";
--            LineBuffer2(1702) <= "00000000";
--            LineBuffer2(1703) <= "00000000";
--            LineBuffer2(1704) <= "00000000";
--            LineBuffer2(1705) <= "00000000";
--            LineBuffer2(1706) <= "00000000";
--            LineBuffer2(1707) <= "00000000";
--            LineBuffer2(1708) <= "00000000";
--            LineBuffer2(1709) <= "00000000";    
--            LineBuffer2(1710) <= "00000000";
--            LineBuffer2(1711) <= "00000000";
--            LineBuffer2(1712) <= "00000000";
--            LineBuffer2(1713) <= "00000000";
--            LineBuffer2(1714) <= "00000000";
--            LineBuffer2(1715) <= "00000000";
--            LineBuffer2(1716) <= "00000000";
--            LineBuffer2(1717) <= "00000000";
--            LineBuffer2(1718) <= "00000000";
--            LineBuffer2(1719) <= "00000000";    
--            LineBuffer2(1720) <= "00000000";
--            LineBuffer2(1721) <= "00000000";
--            LineBuffer2(1722) <= "00000000";
--            LineBuffer2(1723) <= "00000000";
--            LineBuffer2(1724) <= "00000000";
--            LineBuffer2(1725) <= "00000000";
--            LineBuffer2(1726) <= "00000000";
--            LineBuffer2(1727) <= "00000000";
--            LineBuffer2(1728) <= "00000000";
--            LineBuffer2(1729) <= "00000000";    
--            LineBuffer2(1730) <= "00000000";
--            LineBuffer2(1731) <= "00000000";
--            LineBuffer2(1732) <= "00000000";
--            LineBuffer2(1733) <= "00000000";
--            LineBuffer2(1734) <= "00000000";
--            LineBuffer2(1735) <= "00000000";
--            LineBuffer2(1736) <= "00000000";
--            LineBuffer2(1737) <= "00000000";
--            LineBuffer2(1738) <= "00000000";
--            LineBuffer2(1739) <= "00000000";    
--            LineBuffer2(1740) <= "00000000";
--            LineBuffer2(1741) <= "00000000";
--            LineBuffer2(1742) <= "00000000";
--            LineBuffer2(1743) <= "00000000";
--            LineBuffer2(1744) <= "00000000";
--            LineBuffer2(1745) <= "00000000";
--            LineBuffer2(1746) <= "00000000";
--            LineBuffer2(1747) <= "00000000";
--            LineBuffer2(1748) <= "00000000";
--            LineBuffer2(1749) <= "00000000";    
--            LineBuffer2(1750) <= "00000000";
--            LineBuffer2(1751) <= "00000000";
--            LineBuffer2(1752) <= "00000000";
--            LineBuffer2(1753) <= "00000000";
--            LineBuffer2(1754) <= "00000000";
--            LineBuffer2(1755) <= "00000000";
--            LineBuffer2(1756) <= "00000000";
--            LineBuffer2(1757) <= "00000000";
--            LineBuffer2(1758) <= "00000000";
--            LineBuffer2(1759) <= "00000000";    
--            LineBuffer2(1760) <= "00000000";
--            LineBuffer2(1761) <= "00000000";
--            LineBuffer2(1762) <= "00000000";
--            LineBuffer2(1763) <= "00000000";
--            LineBuffer2(1764) <= "00000000";
--            LineBuffer2(1765) <= "00000000";
--            LineBuffer2(1766) <= "00000000";
--            LineBuffer2(1767) <= "00000000";
--            LineBuffer2(1768) <= "00000000";
--            LineBuffer2(1769) <= "00000000";    
--            LineBuffer2(1770) <= "00000000";
--            LineBuffer2(1771) <= "00000000";
--            LineBuffer2(1772) <= "00000000";
--            LineBuffer2(1773) <= "00000000";
--            LineBuffer2(1774) <= "00000000";
--            LineBuffer2(1775) <= "00000000";
--            LineBuffer2(1776) <= "00000000";
--            LineBuffer2(1777) <= "00000000";
--            LineBuffer2(1778) <= "00000000";
--            LineBuffer2(1779) <= "00000000";
--            LineBuffer2(1780) <= "00000000";
--            LineBuffer2(1781) <= "00000000";
--            LineBuffer2(1782) <= "00000000";
--            LineBuffer2(1783) <= "00000000";
--            LineBuffer2(1784) <= "00000000";
--            LineBuffer2(1785) <= "00000000";
--            LineBuffer2(1786) <= "00000000";
--            LineBuffer2(1787) <= "00000000";
--            LineBuffer2(1788) <= "00000000";
--            LineBuffer2(1789) <= "00000000";    
--            LineBuffer2(1790) <= "00000000";
--            LineBuffer2(1791) <= "00000000";
--            LineBuffer2(1792) <= "00000000";
--            LineBuffer2(1793) <= "00000000";
--            LineBuffer2(1794) <= "00000000";
--            LineBuffer2(1795) <= "00000000";
--            LineBuffer2(1796) <= "00000000";
--            LineBuffer2(1797) <= "00000000";
--            LineBuffer2(1798) <= "00000000";
--            LineBuffer2(1799) <= "00000000";    
--            LineBuffer2(1800) <= "00000000";
--            LineBuffer2(1801) <= "00000000";
--            LineBuffer2(1802) <= "00000000";
--            LineBuffer2(1803) <= "00000000";
--            LineBuffer2(1804) <= "00000000";
--            LineBuffer2(1805) <= "00000000";
--            LineBuffer2(1806) <= "00000000";
--            LineBuffer2(1807) <= "00000000";
--            LineBuffer2(1808) <= "00000000";
--            LineBuffer2(1809) <= "00000000";    
--            LineBuffer2(1810) <= "00000000";
--            LineBuffer2(1811) <= "00000000";
--            LineBuffer2(1812) <= "00000000";
--            LineBuffer2(1813) <= "00000000";
--            LineBuffer2(1814) <= "00000000";
--            LineBuffer2(1815) <= "00000000";
--            LineBuffer2(1816) <= "00000000";
--            LineBuffer2(1817) <= "00000000";
--            LineBuffer2(1818) <= "00000000";
--            LineBuffer2(1819) <= "00000000";    
--            LineBuffer2(1820) <= "00000000";
--            LineBuffer2(1821) <= "00000000";
--            LineBuffer2(1822) <= "00000000";
--            LineBuffer2(1823) <= "00000000";
--            LineBuffer2(1824) <= "00000000";
--            LineBuffer2(1825) <= "00000000";
--            LineBuffer2(1826) <= "00000000";
--            LineBuffer2(1827) <= "00000000";
--            LineBuffer2(1828) <= "00000000";
--            LineBuffer2(1829) <= "00000000";    
--            LineBuffer2(1830) <= "00000000";
--            LineBuffer2(1831) <= "00000000";
--            LineBuffer2(1832) <= "00000000";
--            LineBuffer2(1833) <= "00000000";
--            LineBuffer2(1834) <= "00000000";
--            LineBuffer2(1835) <= "00000000";
--            LineBuffer2(1836) <= "00000000";
--            LineBuffer2(1837) <= "00000000";
--            LineBuffer2(1838) <= "00000000";
--            LineBuffer2(1839) <= "00000000";    
--            LineBuffer2(1840) <= "00000000";
--            LineBuffer2(1841) <= "00000000";
--            LineBuffer2(1842) <= "00000000";
--            LineBuffer2(1843) <= "00000000";
--            LineBuffer2(1844) <= "00000000";
--            LineBuffer2(1845) <= "00000000";
--            LineBuffer2(1846) <= "00000000";
--            LineBuffer2(1847) <= "00000000";
--            LineBuffer2(1848) <= "00000000";
--            LineBuffer2(1849) <= "00000000";    
--            LineBuffer2(1850) <= "00000000";
--            LineBuffer2(1851) <= "00000000";
--            LineBuffer2(1852) <= "00000000";
--            LineBuffer2(1853) <= "00000000";
--            LineBuffer2(1854) <= "00000000";
--            LineBuffer2(1855) <= "00000000";
--            LineBuffer2(1856) <= "00000000";
--            LineBuffer2(1857) <= "00000000";
--            LineBuffer2(1858) <= "00000000";
--            LineBuffer2(1859) <= "00000000";    
--            LineBuffer2(1860) <= "00000000";
--            LineBuffer2(1861) <= "00000000";
--            LineBuffer2(1862) <= "00000000";
--            LineBuffer2(1863) <= "00000000";
--            LineBuffer2(1864) <= "00000000";
--            LineBuffer2(1865) <= "00000000";
--            LineBuffer2(1866) <= "00000000";
--            LineBuffer2(1867) <= "00000000";
--            LineBuffer2(1868) <= "00000000";
--            LineBuffer2(1869) <= "00000000";    
--            LineBuffer2(1870) <= "00000000";
--            LineBuffer2(1871) <= "00000000";
--            LineBuffer2(1872) <= "00000000";
--            LineBuffer2(1873) <= "00000000";
--            LineBuffer2(1874) <= "00000000";
--            LineBuffer2(1875) <= "00000000";
--            LineBuffer2(1876) <= "00000000";
--            LineBuffer2(1877) <= "00000000";
--            LineBuffer2(1878) <= "00000000";
--            LineBuffer2(1879) <= "00000000";
--            LineBuffer2(1880) <= "00000000";
--            LineBuffer2(1881) <= "00000000";
--            LineBuffer2(1882) <= "00000000";
--            LineBuffer2(1883) <= "00000000";
--            LineBuffer2(1884) <= "00000000";
--            LineBuffer2(1885) <= "00000000";
--            LineBuffer2(1886) <= "00000000";
--            LineBuffer2(1887) <= "00000000";
--            LineBuffer2(1888) <= "00000000";
--            LineBuffer2(1889) <= "00000000";    
--            LineBuffer2(1890) <= "00000000";
--            LineBuffer2(1891) <= "00000000";
--            LineBuffer2(1892) <= "00000000";
--            LineBuffer2(1893) <= "00000000";
--            LineBuffer2(1894) <= "00000000";
--            LineBuffer2(1895) <= "00000000";
--            LineBuffer2(1896) <= "00000000";
--            LineBuffer2(1897) <= "00000000";
--            LineBuffer2(1898) <= "00000000";
--            LineBuffer2(1899) <= "00000000";    
--            LineBuffer2(1900) <= "00000000";
--            LineBuffer2(1901) <= "00000000";
--            LineBuffer2(1902) <= "00000000";
--            LineBuffer2(1903) <= "00000000";
--            LineBuffer2(1904) <= "00000000";
--            LineBuffer2(1905) <= "00000000";
--            LineBuffer2(1906) <= "00000000";
--            LineBuffer2(1907) <= "00000000";
--            LineBuffer2(1908) <= "00000000";
--            LineBuffer2(1909) <= "00000000";    
--            LineBuffer2(1910) <= "00000000";
--            LineBuffer2(1911) <= "00000000";
--            LineBuffer2(1912) <= "00000000";
--            LineBuffer2(1913) <= "00000000";
--            LineBuffer2(1914) <= "00000000";
--            LineBuffer2(1915) <= "00000000";
--            LineBuffer2(1916) <= "00000000";
--            LineBuffer2(1917) <= "00000000";
--            LineBuffer2(1918) <= "00000000";
--            LineBuffer2(1919) <= "00000000";	
			
			
			
			
			
						
				else
	        LineBuffer0(0) <= shiftin;	
			LineBuffer0(1) <= LineBuffer0(0);
			LineBuffer0(2) <= LineBuffer0(1);
			LineBuffer0(3) <= LineBuffer0(2);
			LineBuffer0(4) <= LineBuffer0(3);
			LineBuffer0(5) <= LineBuffer0(4);
			LineBuffer0(6) <= LineBuffer0(5);
			LineBuffer0(7) <= LineBuffer0(6);
			LineBuffer0(8) <= LineBuffer0(7);
			LineBuffer0(9) <= LineBuffer0(8);	
			LineBuffer0(10) <= LineBuffer0(9);
			LineBuffer0(11) <= LineBuffer0(10);
			LineBuffer0(12) <= LineBuffer0(11);
			LineBuffer0(13) <= LineBuffer0(12);
			LineBuffer0(14) <= LineBuffer0(13);
			LineBuffer0(15) <= LineBuffer0(14);
			LineBuffer0(16) <= LineBuffer0(15);
			LineBuffer0(17) <= LineBuffer0(16);
			LineBuffer0(18) <= LineBuffer0(17);
			LineBuffer0(19) <= LineBuffer0(18);	
			LineBuffer0(20) <= LineBuffer0(19);
			LineBuffer0(21) <= LineBuffer0(20);
			LineBuffer0(22) <= LineBuffer0(21);
			LineBuffer0(23) <= LineBuffer0(22);
			LineBuffer0(24) <= LineBuffer0(23);
			LineBuffer0(25) <= LineBuffer0(24);
			LineBuffer0(26) <= LineBuffer0(25);
			LineBuffer0(27) <= LineBuffer0(26);
			LineBuffer0(28) <= LineBuffer0(27);
			LineBuffer0(29) <= LineBuffer0(28);	
			LineBuffer0(30) <= LineBuffer0(29);
			LineBuffer0(31) <= LineBuffer0(30);
			LineBuffer0(32) <= LineBuffer0(31);
			LineBuffer0(33) <= LineBuffer0(32);
			LineBuffer0(34) <= LineBuffer0(33);
			LineBuffer0(35) <= LineBuffer0(34);
			LineBuffer0(36) <= LineBuffer0(35);
			LineBuffer0(37) <= LineBuffer0(36);
			LineBuffer0(38) <= LineBuffer0(37);
			LineBuffer0(39) <= LineBuffer0(38);	
			LineBuffer0(40) <= LineBuffer0(39);
			LineBuffer0(41) <= LineBuffer0(40);
			LineBuffer0(42) <= LineBuffer0(41);
			LineBuffer0(43) <= LineBuffer0(42);
			LineBuffer0(44) <= LineBuffer0(43);
			LineBuffer0(45) <= LineBuffer0(44);
			LineBuffer0(46) <= LineBuffer0(45);
			LineBuffer0(47) <= LineBuffer0(46);
			LineBuffer0(48) <= LineBuffer0(47);
			LineBuffer0(49) <= LineBuffer0(48);	
			LineBuffer0(50) <= LineBuffer0(49);
			LineBuffer0(51) <= LineBuffer0(50);
			LineBuffer0(52) <= LineBuffer0(51);
			LineBuffer0(53) <= LineBuffer0(52);
			LineBuffer0(54) <= LineBuffer0(53);
			LineBuffer0(55) <= LineBuffer0(54);
			LineBuffer0(56) <= LineBuffer0(55);
			LineBuffer0(57) <= LineBuffer0(56);
			LineBuffer0(58) <= LineBuffer0(57);
			LineBuffer0(59) <= LineBuffer0(58);	
			LineBuffer0(60) <= LineBuffer0(59);
			LineBuffer0(61) <= LineBuffer0(60);
			LineBuffer0(62) <= LineBuffer0(61);
			LineBuffer0(63) <= LineBuffer0(62);
			LineBuffer0(64) <= LineBuffer0(63);
			LineBuffer0(65) <= LineBuffer0(64);
			LineBuffer0(66) <= LineBuffer0(65);
			LineBuffer0(67) <= LineBuffer0(66);
			LineBuffer0(68) <= LineBuffer0(67);
			LineBuffer0(69) <= LineBuffer0(68);	
			LineBuffer0(70) <= LineBuffer0(69);
			LineBuffer0(71) <= LineBuffer0(70);
			LineBuffer0(72) <= LineBuffer0(71);
			LineBuffer0(73) <= LineBuffer0(72);
			LineBuffer0(74) <= LineBuffer0(73);
			LineBuffer0(75) <= LineBuffer0(74);
			LineBuffer0(76) <= LineBuffer0(75);
			LineBuffer0(77) <= LineBuffer0(76);
			LineBuffer0(78) <= LineBuffer0(77);
			LineBuffer0(79) <= LineBuffer0(78);	
			LineBuffer0(80) <= LineBuffer0(79);
			LineBuffer0(81) <= LineBuffer0(80);
			LineBuffer0(82) <= LineBuffer0(81);
			LineBuffer0(83) <= LineBuffer0(82);
			LineBuffer0(84) <= LineBuffer0(83);
			LineBuffer0(85) <= LineBuffer0(84);
			LineBuffer0(86) <= LineBuffer0(85);
			LineBuffer0(87) <= LineBuffer0(86);
			LineBuffer0(88) <= LineBuffer0(87);
			LineBuffer0(89) <= LineBuffer0(88);	
			LineBuffer0(90) <= LineBuffer0(89);
			LineBuffer0(91) <= LineBuffer0(90);
			LineBuffer0(92) <= LineBuffer0(91);
			LineBuffer0(93) <= LineBuffer0(92);
			LineBuffer0(94) <= LineBuffer0(93);
			LineBuffer0(95) <= LineBuffer0(94);
			LineBuffer0(96) <= LineBuffer0(95);
			LineBuffer0(97) <= LineBuffer0(96);
			LineBuffer0(98) <= LineBuffer0(97);
			LineBuffer0(99) <= LineBuffer0(98);	
			LineBuffer0(100) <= LineBuffer0(99);
			LineBuffer0(101) <= LineBuffer0(100);
			LineBuffer0(102) <= LineBuffer0(101);
			LineBuffer0(103) <= LineBuffer0(102);
			LineBuffer0(104) <= LineBuffer0(103);
			LineBuffer0(105) <= LineBuffer0(104);
			LineBuffer0(106) <= LineBuffer0(105);
			LineBuffer0(107) <= LineBuffer0(106);
			LineBuffer0(108) <= LineBuffer0(107);
			LineBuffer0(109) <= LineBuffer0(108);	
			LineBuffer0(110) <= LineBuffer0(109);
			LineBuffer0(111) <= LineBuffer0(110);
			LineBuffer0(112) <= LineBuffer0(111);
			LineBuffer0(113) <= LineBuffer0(112);
			LineBuffer0(114) <= LineBuffer0(113);
			LineBuffer0(115) <= LineBuffer0(114);
			LineBuffer0(116) <= LineBuffer0(115);
			LineBuffer0(117) <= LineBuffer0(116);
			LineBuffer0(118) <= LineBuffer0(117);
			LineBuffer0(119) <= LineBuffer0(118);	
			LineBuffer0(120) <= LineBuffer0(119);
			LineBuffer0(121) <= LineBuffer0(120);
			LineBuffer0(122) <= LineBuffer0(121);
			LineBuffer0(123) <= LineBuffer0(122);
			LineBuffer0(124) <= LineBuffer0(123);
			LineBuffer0(125) <= LineBuffer0(124);
			LineBuffer0(126) <= LineBuffer0(125);
			LineBuffer0(127) <= LineBuffer0(126);
			LineBuffer0(128) <= LineBuffer0(127);
			LineBuffer0(129) <= LineBuffer0(128);	
			LineBuffer0(130) <= LineBuffer0(129);
			LineBuffer0(131) <= LineBuffer0(130);
			LineBuffer0(132) <= LineBuffer0(131);
			LineBuffer0(133) <= LineBuffer0(132);
			LineBuffer0(134) <= LineBuffer0(133);
			LineBuffer0(135) <= LineBuffer0(134);
			LineBuffer0(136) <= LineBuffer0(135);
			LineBuffer0(137) <= LineBuffer0(136);
			LineBuffer0(138) <= LineBuffer0(137);
			LineBuffer0(139) <= LineBuffer0(138);	
			LineBuffer0(140) <= LineBuffer0(139);
			LineBuffer0(141) <= LineBuffer0(140);
			LineBuffer0(142) <= LineBuffer0(141);
			LineBuffer0(143) <= LineBuffer0(142);
			LineBuffer0(144) <= LineBuffer0(143);
			LineBuffer0(145) <= LineBuffer0(144);
			LineBuffer0(146) <= LineBuffer0(145);
			LineBuffer0(147) <= LineBuffer0(146);
			LineBuffer0(148) <= LineBuffer0(147);
			LineBuffer0(149) <= LineBuffer0(148);	
			LineBuffer0(150) <= LineBuffer0(149);
			LineBuffer0(151) <= LineBuffer0(150);
			LineBuffer0(152) <= LineBuffer0(151);
			LineBuffer0(153) <= LineBuffer0(152);
			LineBuffer0(154) <= LineBuffer0(153);
			LineBuffer0(155) <= LineBuffer0(154);
			LineBuffer0(156) <= LineBuffer0(155);
			LineBuffer0(157) <= LineBuffer0(156);
			LineBuffer0(158) <= LineBuffer0(157);
			LineBuffer0(159) <= LineBuffer0(158);	
			LineBuffer0(160) <= LineBuffer0(159);
			LineBuffer0(161) <= LineBuffer0(160);
			LineBuffer0(162) <= LineBuffer0(161);
			LineBuffer0(163) <= LineBuffer0(162);
			LineBuffer0(164) <= LineBuffer0(163);
			LineBuffer0(165) <= LineBuffer0(164);
			LineBuffer0(166) <= LineBuffer0(165);
			LineBuffer0(167) <= LineBuffer0(166);
			LineBuffer0(168) <= LineBuffer0(167);
			LineBuffer0(169) <= LineBuffer0(168);	
			LineBuffer0(170) <= LineBuffer0(169);
			LineBuffer0(171) <= LineBuffer0(170);
			LineBuffer0(172) <= LineBuffer0(171);
			LineBuffer0(173) <= LineBuffer0(172);
			LineBuffer0(174) <= LineBuffer0(173);
			LineBuffer0(175) <= LineBuffer0(174);
			LineBuffer0(176) <= LineBuffer0(175);
			LineBuffer0(177) <= LineBuffer0(176);
			LineBuffer0(178) <= LineBuffer0(177);
			LineBuffer0(179) <= LineBuffer0(178);	
			LineBuffer0(180) <= LineBuffer0(179);
			LineBuffer0(181) <= LineBuffer0(180);
			LineBuffer0(182) <= LineBuffer0(181);
			LineBuffer0(183) <= LineBuffer0(182);
			LineBuffer0(184) <= LineBuffer0(183);
			LineBuffer0(185) <= LineBuffer0(184);
			LineBuffer0(186) <= LineBuffer0(185);
			LineBuffer0(187) <= LineBuffer0(186);
			LineBuffer0(188) <= LineBuffer0(187);
			LineBuffer0(189) <= LineBuffer0(188);	
			LineBuffer0(190) <= LineBuffer0(189);
			LineBuffer0(191) <= LineBuffer0(190);
			LineBuffer0(192) <= LineBuffer0(191);
			LineBuffer0(193) <= LineBuffer0(192);
			LineBuffer0(194) <= LineBuffer0(193);
			LineBuffer0(195) <= LineBuffer0(194);
			LineBuffer0(196) <= LineBuffer0(195);
			LineBuffer0(197) <= LineBuffer0(196);
			LineBuffer0(198) <= LineBuffer0(197);
			LineBuffer0(199) <= LineBuffer0(198);
			LineBuffer0(200) <= LineBuffer0(199);
			LineBuffer0(201) <= LineBuffer0(200);
			LineBuffer0(202) <= LineBuffer0(201);
			LineBuffer0(203) <= LineBuffer0(202);
			LineBuffer0(204) <= LineBuffer0(203);
			LineBuffer0(205) <= LineBuffer0(204);
			LineBuffer0(206) <= LineBuffer0(205);
			LineBuffer0(207) <= LineBuffer0(206);
			LineBuffer0(208) <= LineBuffer0(207);
			LineBuffer0(209) <= LineBuffer0(208);	
			LineBuffer0(210) <= LineBuffer0(209);
			LineBuffer0(211) <= LineBuffer0(210);
			LineBuffer0(212) <= LineBuffer0(211);
			LineBuffer0(213) <= LineBuffer0(212);
			LineBuffer0(214) <= LineBuffer0(213);
			LineBuffer0(215) <= LineBuffer0(214);
			LineBuffer0(216) <= LineBuffer0(215);
			LineBuffer0(217) <= LineBuffer0(216);
			LineBuffer0(218) <= LineBuffer0(217);
			LineBuffer0(219) <= LineBuffer0(218);	
			LineBuffer0(220) <= LineBuffer0(219);
			LineBuffer0(221) <= LineBuffer0(220);
			LineBuffer0(222) <= LineBuffer0(221);
			LineBuffer0(223) <= LineBuffer0(222);
			LineBuffer0(224) <= LineBuffer0(223);
			LineBuffer0(225) <= LineBuffer0(224);
			LineBuffer0(226) <= LineBuffer0(225);
			LineBuffer0(227) <= LineBuffer0(226);
			LineBuffer0(228) <= LineBuffer0(227);
			LineBuffer0(229) <= LineBuffer0(228);	
			LineBuffer0(230) <= LineBuffer0(229);
			LineBuffer0(231) <= LineBuffer0(230);
			LineBuffer0(232) <= LineBuffer0(231);
			LineBuffer0(233) <= LineBuffer0(232);
			LineBuffer0(234) <= LineBuffer0(233);
			LineBuffer0(235) <= LineBuffer0(234);
			LineBuffer0(236) <= LineBuffer0(235);
			LineBuffer0(237) <= LineBuffer0(236);
			LineBuffer0(238) <= LineBuffer0(237);
			LineBuffer0(239) <= LineBuffer0(238);	
			LineBuffer0(240) <= LineBuffer0(239);
			LineBuffer0(241) <= LineBuffer0(240);
			LineBuffer0(242) <= LineBuffer0(241);
			LineBuffer0(243) <= LineBuffer0(242);
			LineBuffer0(244) <= LineBuffer0(243);
			LineBuffer0(245) <= LineBuffer0(244);
			LineBuffer0(246) <= LineBuffer0(245);
			LineBuffer0(247) <= LineBuffer0(246);
			LineBuffer0(248) <= LineBuffer0(247);
			LineBuffer0(249) <= LineBuffer0(248);	
			LineBuffer0(250) <= LineBuffer0(249);
			LineBuffer0(251) <= LineBuffer0(250);
			LineBuffer0(252) <= LineBuffer0(251);
			LineBuffer0(253) <= LineBuffer0(252);
			LineBuffer0(254) <= LineBuffer0(253);
			LineBuffer0(255) <= LineBuffer0(254);
			LineBuffer0(256) <= LineBuffer0(255);
			LineBuffer0(257) <= LineBuffer0(256);
			LineBuffer0(258) <= LineBuffer0(257);
			LineBuffer0(259) <= LineBuffer0(258);	
			LineBuffer0(260) <= LineBuffer0(259);
			LineBuffer0(261) <= LineBuffer0(260);
			LineBuffer0(262) <= LineBuffer0(261);
			LineBuffer0(263) <= LineBuffer0(262);
			LineBuffer0(264) <= LineBuffer0(263);
			LineBuffer0(265) <= LineBuffer0(264);
			LineBuffer0(266) <= LineBuffer0(265);
			LineBuffer0(267) <= LineBuffer0(266);
			LineBuffer0(268) <= LineBuffer0(267);
			LineBuffer0(269) <= LineBuffer0(268);	
			LineBuffer0(270) <= LineBuffer0(269);
			LineBuffer0(271) <= LineBuffer0(270);
			LineBuffer0(272) <= LineBuffer0(271);
			LineBuffer0(273) <= LineBuffer0(272);
			LineBuffer0(274) <= LineBuffer0(273);
			LineBuffer0(275) <= LineBuffer0(274);
			LineBuffer0(276) <= LineBuffer0(275);
			LineBuffer0(277) <= LineBuffer0(276);
			LineBuffer0(278) <= LineBuffer0(277);
			LineBuffer0(279) <= LineBuffer0(278);	
			LineBuffer0(280) <= LineBuffer0(279);
			LineBuffer0(281) <= LineBuffer0(280);
			LineBuffer0(282) <= LineBuffer0(281);
			LineBuffer0(283) <= LineBuffer0(282);
			LineBuffer0(284) <= LineBuffer0(283);
			LineBuffer0(285) <= LineBuffer0(284);
			LineBuffer0(286) <= LineBuffer0(285);
			LineBuffer0(287) <= LineBuffer0(286);
			LineBuffer0(288) <= LineBuffer0(287);
			LineBuffer0(289) <= LineBuffer0(288);	
			LineBuffer0(290) <= LineBuffer0(289);
			LineBuffer0(291) <= LineBuffer0(290);
			LineBuffer0(292) <= LineBuffer0(291);
			LineBuffer0(293) <= LineBuffer0(292);
			LineBuffer0(294) <= LineBuffer0(293);
			LineBuffer0(295) <= LineBuffer0(294);
			LineBuffer0(296) <= LineBuffer0(295);
			LineBuffer0(297) <= LineBuffer0(296);
			LineBuffer0(298) <= LineBuffer0(297);
			LineBuffer0(299) <= LineBuffer0(298);	
			LineBuffer0(300) <= LineBuffer0(299);	
			LineBuffer0(301) <= LineBuffer0(300);
			LineBuffer0(302) <= LineBuffer0(301);
			LineBuffer0(303) <= LineBuffer0(302);
			LineBuffer0(304) <= LineBuffer0(303);
			LineBuffer0(305) <= LineBuffer0(304);
			LineBuffer0(306) <= LineBuffer0(305);
			LineBuffer0(307) <= LineBuffer0(306);
			LineBuffer0(308) <= LineBuffer0(307);
			LineBuffer0(309) <= LineBuffer0(308);	
			LineBuffer0(310) <= LineBuffer0(309);
			LineBuffer0(311) <= LineBuffer0(310);
			LineBuffer0(312) <= LineBuffer0(311);
			LineBuffer0(313) <= LineBuffer0(312);
			LineBuffer0(314) <= LineBuffer0(313);
			LineBuffer0(315) <= LineBuffer0(314);
			LineBuffer0(316) <= LineBuffer0(315);
			LineBuffer0(317) <= LineBuffer0(316);
			LineBuffer0(318) <= LineBuffer0(317);
			LineBuffer0(319) <= LineBuffer0(318);	
			LineBuffer0(320) <= LineBuffer0(319);
			LineBuffer0(321) <= LineBuffer0(320);
			LineBuffer0(322) <= LineBuffer0(321);
			LineBuffer0(323) <= LineBuffer0(322);
			LineBuffer0(324) <= LineBuffer0(323);
			LineBuffer0(325) <= LineBuffer0(324);
			LineBuffer0(326) <= LineBuffer0(325);
			LineBuffer0(327) <= LineBuffer0(326);
			LineBuffer0(328) <= LineBuffer0(327);
			LineBuffer0(329) <= LineBuffer0(328);	
			LineBuffer0(330) <= LineBuffer0(329);
			LineBuffer0(331) <= LineBuffer0(330);
			LineBuffer0(332) <= LineBuffer0(331);
			LineBuffer0(333) <= LineBuffer0(332);
			LineBuffer0(334) <= LineBuffer0(333);
			LineBuffer0(335) <= LineBuffer0(334);
			LineBuffer0(336) <= LineBuffer0(335);
			LineBuffer0(337) <= LineBuffer0(336);
			LineBuffer0(338) <= LineBuffer0(337);
			LineBuffer0(339) <= LineBuffer0(338);	
			LineBuffer0(340) <= LineBuffer0(339);
			LineBuffer0(341) <= LineBuffer0(340);
			LineBuffer0(342) <= LineBuffer0(341);
			LineBuffer0(343) <= LineBuffer0(342);
			LineBuffer0(344) <= LineBuffer0(343);
			LineBuffer0(345) <= LineBuffer0(344);
			LineBuffer0(346) <= LineBuffer0(345);
			LineBuffer0(347) <= LineBuffer0(346);
			LineBuffer0(348) <= LineBuffer0(347);
			LineBuffer0(349) <= LineBuffer0(348);	
			LineBuffer0(350) <= LineBuffer0(349);
			LineBuffer0(351) <= LineBuffer0(350);
			LineBuffer0(352) <= LineBuffer0(351);
			LineBuffer0(353) <= LineBuffer0(352);
			LineBuffer0(354) <= LineBuffer0(353);
			LineBuffer0(355) <= LineBuffer0(354);
			LineBuffer0(356) <= LineBuffer0(355);
			LineBuffer0(357) <= LineBuffer0(356);
			LineBuffer0(358) <= LineBuffer0(357);
			LineBuffer0(359) <= LineBuffer0(358);	
			LineBuffer0(360) <= LineBuffer0(359);
			LineBuffer0(361) <= LineBuffer0(360);
			LineBuffer0(362) <= LineBuffer0(361);
			LineBuffer0(363) <= LineBuffer0(362);
			LineBuffer0(364) <= LineBuffer0(363);
			LineBuffer0(365) <= LineBuffer0(364);
			LineBuffer0(366) <= LineBuffer0(365);
			LineBuffer0(367) <= LineBuffer0(366);
			LineBuffer0(368) <= LineBuffer0(367);
			LineBuffer0(369) <= LineBuffer0(368);	
			LineBuffer0(370) <= LineBuffer0(369);
			LineBuffer0(371) <= LineBuffer0(370);
			LineBuffer0(372) <= LineBuffer0(371);
			LineBuffer0(373) <= LineBuffer0(372);
			LineBuffer0(374) <= LineBuffer0(373);
			LineBuffer0(375) <= LineBuffer0(374);
			LineBuffer0(376) <= LineBuffer0(375);
			LineBuffer0(377) <= LineBuffer0(376);
			LineBuffer0(378) <= LineBuffer0(377);
			LineBuffer0(379) <= LineBuffer0(378);	
			LineBuffer0(380) <= LineBuffer0(379);
			LineBuffer0(381) <= LineBuffer0(380);
			LineBuffer0(382) <= LineBuffer0(381);
			LineBuffer0(383) <= LineBuffer0(382);
			LineBuffer0(384) <= LineBuffer0(383);
			LineBuffer0(385) <= LineBuffer0(384);
			LineBuffer0(386) <= LineBuffer0(385);
			LineBuffer0(387) <= LineBuffer0(386);
			LineBuffer0(388) <= LineBuffer0(387);
			LineBuffer0(389) <= LineBuffer0(388);	
			LineBuffer0(390) <= LineBuffer0(389);
			LineBuffer0(391) <= LineBuffer0(390);
			LineBuffer0(392) <= LineBuffer0(391);
			LineBuffer0(393) <= LineBuffer0(392);
			LineBuffer0(394) <= LineBuffer0(393);
			LineBuffer0(395) <= LineBuffer0(394);
			LineBuffer0(396) <= LineBuffer0(395);
			LineBuffer0(397) <= LineBuffer0(396);
			LineBuffer0(398) <= LineBuffer0(397);
			LineBuffer0(399) <= LineBuffer0(398);
			LineBuffer0(400) <= LineBuffer0(399);	
			LineBuffer0(401) <= LineBuffer0(400);
			LineBuffer0(402) <= LineBuffer0(401);
			LineBuffer0(403) <= LineBuffer0(402);
			LineBuffer0(404) <= LineBuffer0(403);
			LineBuffer0(405) <= LineBuffer0(404);
			LineBuffer0(406) <= LineBuffer0(405);
			LineBuffer0(407) <= LineBuffer0(406);
			LineBuffer0(408) <= LineBuffer0(407);
			LineBuffer0(409) <= LineBuffer0(408);	
			LineBuffer0(410) <= LineBuffer0(409);
			LineBuffer0(411) <= LineBuffer0(410);
			LineBuffer0(412) <= LineBuffer0(411);
			LineBuffer0(413) <= LineBuffer0(412);
			LineBuffer0(414) <= LineBuffer0(413);
			LineBuffer0(415) <= LineBuffer0(414);
			LineBuffer0(416) <= LineBuffer0(415);
			LineBuffer0(417) <= LineBuffer0(416);
			LineBuffer0(418) <= LineBuffer0(417);
			LineBuffer0(419) <= LineBuffer0(418);	
			LineBuffer0(420) <= LineBuffer0(419);
			LineBuffer0(421) <= LineBuffer0(420);
			LineBuffer0(422) <= LineBuffer0(421);
			LineBuffer0(423) <= LineBuffer0(422);
			LineBuffer0(424) <= LineBuffer0(423);
			LineBuffer0(425) <= LineBuffer0(424);
			LineBuffer0(426) <= LineBuffer0(425);
			LineBuffer0(427) <= LineBuffer0(426);
			LineBuffer0(428) <= LineBuffer0(427);
			LineBuffer0(429) <= LineBuffer0(428);	
			LineBuffer0(430) <= LineBuffer0(429);
			LineBuffer0(431) <= LineBuffer0(430);
			LineBuffer0(432) <= LineBuffer0(431);
			LineBuffer0(433) <= LineBuffer0(432);
			LineBuffer0(434) <= LineBuffer0(433);
			LineBuffer0(435) <= LineBuffer0(434);
			LineBuffer0(436) <= LineBuffer0(435);
			LineBuffer0(437) <= LineBuffer0(436);
			LineBuffer0(438) <= LineBuffer0(437);
			LineBuffer0(439) <= LineBuffer0(438);	
			LineBuffer0(440) <= LineBuffer0(439);
			LineBuffer0(441) <= LineBuffer0(440);
			LineBuffer0(442) <= LineBuffer0(441);
			LineBuffer0(443) <= LineBuffer0(442);
			LineBuffer0(444) <= LineBuffer0(443);
			LineBuffer0(445) <= LineBuffer0(444);
			LineBuffer0(446) <= LineBuffer0(445);
			LineBuffer0(447) <= LineBuffer0(446);
			LineBuffer0(448) <= LineBuffer0(447);
			LineBuffer0(449) <= LineBuffer0(448);	
			LineBuffer0(450) <= LineBuffer0(449);
			LineBuffer0(451) <= LineBuffer0(450);
			LineBuffer0(452) <= LineBuffer0(451);
			LineBuffer0(453) <= LineBuffer0(452);
			LineBuffer0(454) <= LineBuffer0(453);
			LineBuffer0(455) <= LineBuffer0(454);
			LineBuffer0(456) <= LineBuffer0(455);
			LineBuffer0(457) <= LineBuffer0(456);
			LineBuffer0(458) <= LineBuffer0(457);
			LineBuffer0(459) <= LineBuffer0(458);	
			LineBuffer0(460) <= LineBuffer0(459);
			LineBuffer0(461) <= LineBuffer0(460);
			LineBuffer0(462) <= LineBuffer0(461);
			LineBuffer0(463) <= LineBuffer0(462);
			LineBuffer0(464) <= LineBuffer0(463);
			LineBuffer0(465) <= LineBuffer0(464);
			LineBuffer0(466) <= LineBuffer0(465);
			LineBuffer0(467) <= LineBuffer0(466);
			LineBuffer0(468) <= LineBuffer0(467);
			LineBuffer0(469) <= LineBuffer0(468);	
			LineBuffer0(470) <= LineBuffer0(469);
			LineBuffer0(471) <= LineBuffer0(470);
			LineBuffer0(472) <= LineBuffer0(471);
			LineBuffer0(473) <= LineBuffer0(472);
			LineBuffer0(474) <= LineBuffer0(473);
			LineBuffer0(475) <= LineBuffer0(474);
			LineBuffer0(476) <= LineBuffer0(475);
			LineBuffer0(477) <= LineBuffer0(476);
			LineBuffer0(478) <= LineBuffer0(477);
			LineBuffer0(479) <= LineBuffer0(478);	
			LineBuffer0(480) <= LineBuffer0(479);
			LineBuffer0(481) <= LineBuffer0(480);
			LineBuffer0(482) <= LineBuffer0(481);
			LineBuffer0(483) <= LineBuffer0(482);
			LineBuffer0(484) <= LineBuffer0(483);
			LineBuffer0(485) <= LineBuffer0(484);
			LineBuffer0(486) <= LineBuffer0(485);
			LineBuffer0(487) <= LineBuffer0(486);
			LineBuffer0(488) <= LineBuffer0(487);
			LineBuffer0(489) <= LineBuffer0(488);	
			LineBuffer0(490) <= LineBuffer0(489);
			LineBuffer0(491) <= LineBuffer0(490);
			LineBuffer0(492) <= LineBuffer0(491);
			LineBuffer0(493) <= LineBuffer0(492);
			LineBuffer0(494) <= LineBuffer0(493);
			LineBuffer0(495) <= LineBuffer0(494);
			LineBuffer0(496) <= LineBuffer0(495);
			LineBuffer0(497) <= LineBuffer0(496);
			LineBuffer0(498) <= LineBuffer0(497);
			LineBuffer0(499) <= LineBuffer0(498);	
			LineBuffer0(500) <= LineBuffer0(499);	
			LineBuffer0(501) <= LineBuffer0(500);
			LineBuffer0(502) <= LineBuffer0(501);
			LineBuffer0(503) <= LineBuffer0(502);
			LineBuffer0(504) <= LineBuffer0(503);
			LineBuffer0(505) <= LineBuffer0(504);
			LineBuffer0(506) <= LineBuffer0(505);
			LineBuffer0(507) <= LineBuffer0(506);
			LineBuffer0(508) <= LineBuffer0(507);
			LineBuffer0(509) <= LineBuffer0(508);	
			LineBuffer0(510) <= LineBuffer0(509);
			LineBuffer0(511) <= LineBuffer0(510);
			LineBuffer0(512) <= LineBuffer0(511);
			LineBuffer0(513) <= LineBuffer0(512);
			LineBuffer0(514) <= LineBuffer0(513);
			LineBuffer0(515) <= LineBuffer0(514);
			LineBuffer0(516) <= LineBuffer0(515);
			LineBuffer0(517) <= LineBuffer0(516);
			LineBuffer0(518) <= LineBuffer0(517);
			LineBuffer0(519) <= LineBuffer0(518);	
			LineBuffer0(520) <= LineBuffer0(519);
			LineBuffer0(521) <= LineBuffer0(520);
			LineBuffer0(522) <= LineBuffer0(521);
			LineBuffer0(523) <= LineBuffer0(522);
			LineBuffer0(524) <= LineBuffer0(523);
			LineBuffer0(525) <= LineBuffer0(524);
			LineBuffer0(526) <= LineBuffer0(525);
			LineBuffer0(527) <= LineBuffer0(526);
			LineBuffer0(528) <= LineBuffer0(527);
			LineBuffer0(529) <= LineBuffer0(528);	
			LineBuffer0(530) <= LineBuffer0(529);
			LineBuffer0(531) <= LineBuffer0(530);
			LineBuffer0(532) <= LineBuffer0(531);
			LineBuffer0(533) <= LineBuffer0(532);
			LineBuffer0(534) <= LineBuffer0(533);
			LineBuffer0(535) <= LineBuffer0(534);
			LineBuffer0(536) <= LineBuffer0(535);
			LineBuffer0(537) <= LineBuffer0(536);
			LineBuffer0(538) <= LineBuffer0(537);
			LineBuffer0(539) <= LineBuffer0(538);	
			LineBuffer0(540) <= LineBuffer0(539);
			LineBuffer0(541) <= LineBuffer0(540);
			LineBuffer0(542) <= LineBuffer0(541);
			LineBuffer0(543) <= LineBuffer0(542);
			LineBuffer0(544) <= LineBuffer0(543);
			LineBuffer0(545) <= LineBuffer0(544);
			LineBuffer0(546) <= LineBuffer0(545);
			LineBuffer0(547) <= LineBuffer0(546);
			LineBuffer0(548) <= LineBuffer0(547);
			LineBuffer0(549) <= LineBuffer0(548);	
			LineBuffer0(550) <= LineBuffer0(549);
			LineBuffer0(551) <= LineBuffer0(550);
			LineBuffer0(552) <= LineBuffer0(551);
			LineBuffer0(553) <= LineBuffer0(552);
			LineBuffer0(554) <= LineBuffer0(553);
			LineBuffer0(555) <= LineBuffer0(554);
			LineBuffer0(556) <= LineBuffer0(555);
			LineBuffer0(557) <= LineBuffer0(556);
			LineBuffer0(558) <= LineBuffer0(557);
			LineBuffer0(559) <= LineBuffer0(558);	
			LineBuffer0(560) <= LineBuffer0(559);
			LineBuffer0(561) <= LineBuffer0(560);
			LineBuffer0(562) <= LineBuffer0(561);
			LineBuffer0(563) <= LineBuffer0(562);
			LineBuffer0(564) <= LineBuffer0(563);
			LineBuffer0(565) <= LineBuffer0(564);
			LineBuffer0(566) <= LineBuffer0(565);
			LineBuffer0(567) <= LineBuffer0(566);
			LineBuffer0(568) <= LineBuffer0(567);
			LineBuffer0(569) <= LineBuffer0(568);	
			LineBuffer0(570) <= LineBuffer0(569);
			LineBuffer0(571) <= LineBuffer0(570);
			LineBuffer0(572) <= LineBuffer0(571);
			LineBuffer0(573) <= LineBuffer0(572);
			LineBuffer0(574) <= LineBuffer0(573);
			LineBuffer0(575) <= LineBuffer0(574);
			LineBuffer0(576) <= LineBuffer0(575);
			LineBuffer0(577) <= LineBuffer0(576);
			LineBuffer0(578) <= LineBuffer0(577);
			LineBuffer0(579) <= LineBuffer0(578);	
			LineBuffer0(580) <= LineBuffer0(579);
			LineBuffer0(581) <= LineBuffer0(580);
			LineBuffer0(582) <= LineBuffer0(581);
			LineBuffer0(583) <= LineBuffer0(582);
			LineBuffer0(584) <= LineBuffer0(583);
			LineBuffer0(585) <= LineBuffer0(584);
			LineBuffer0(586) <= LineBuffer0(585);
			LineBuffer0(587) <= LineBuffer0(586);
			LineBuffer0(588) <= LineBuffer0(587);
			LineBuffer0(589) <= LineBuffer0(588);	
			LineBuffer0(590) <= LineBuffer0(589);
			LineBuffer0(591) <= LineBuffer0(590);
			LineBuffer0(592) <= LineBuffer0(591);
			LineBuffer0(593) <= LineBuffer0(592);
			LineBuffer0(594) <= LineBuffer0(593);
			LineBuffer0(595) <= LineBuffer0(594);
			LineBuffer0(596) <= LineBuffer0(595);
			LineBuffer0(597) <= LineBuffer0(596);
			LineBuffer0(598) <= LineBuffer0(597);
			LineBuffer0(599) <= LineBuffer0(598);	
			LineBuffer0(600) <= LineBuffer0(599);	
			LineBuffer0(601) <= LineBuffer0(600);
			LineBuffer0(602) <= LineBuffer0(601);
			LineBuffer0(603) <= LineBuffer0(602);
			LineBuffer0(604) <= LineBuffer0(603);
			LineBuffer0(605) <= LineBuffer0(604);
			LineBuffer0(606) <= LineBuffer0(605);
			LineBuffer0(607) <= LineBuffer0(606);
			LineBuffer0(608) <= LineBuffer0(607);
			LineBuffer0(609) <= LineBuffer0(608);	
			LineBuffer0(610) <= LineBuffer0(609);
			LineBuffer0(611) <= LineBuffer0(610);
			LineBuffer0(612) <= LineBuffer0(611);
			LineBuffer0(613) <= LineBuffer0(612);
			LineBuffer0(614) <= LineBuffer0(613);
			LineBuffer0(615) <= LineBuffer0(614);
			LineBuffer0(616) <= LineBuffer0(615);
			LineBuffer0(617) <= LineBuffer0(616);
			LineBuffer0(618) <= LineBuffer0(617);
			LineBuffer0(619) <= LineBuffer0(618);	
			LineBuffer0(620) <= LineBuffer0(619);
			LineBuffer0(621) <= LineBuffer0(620);
			LineBuffer0(622) <= LineBuffer0(621);
			LineBuffer0(623) <= LineBuffer0(622);
			LineBuffer0(624) <= LineBuffer0(623);
			LineBuffer0(625) <= LineBuffer0(624);
			LineBuffer0(626) <= LineBuffer0(625);
			LineBuffer0(627) <= LineBuffer0(626);
			LineBuffer0(628) <= LineBuffer0(627);
			LineBuffer0(629) <= LineBuffer0(628);	
			LineBuffer0(630) <= LineBuffer0(629);
			LineBuffer0(631) <= LineBuffer0(630);
			LineBuffer0(632) <= LineBuffer0(631);
			LineBuffer0(633) <= LineBuffer0(632);
			LineBuffer0(634) <= LineBuffer0(633);
			LineBuffer0(635) <= LineBuffer0(634);
			LineBuffer0(636) <= LineBuffer0(635);
			LineBuffer0(637) <= LineBuffer0(636);
			LineBuffer0(638) <= LineBuffer0(637);
			LineBuffer0(639) <= LineBuffer0(638);
			LineBuffer0(640) <= LineBuffer0(639);
            LineBuffer0(641) <= LineBuffer0(640);
            LineBuffer0(642) <= LineBuffer0(641);
            LineBuffer0(643) <= LineBuffer0(642);
            LineBuffer0(644) <= LineBuffer0(643);
            LineBuffer0(645) <= LineBuffer0(644);
            LineBuffer0(646) <= LineBuffer0(645);
            LineBuffer0(647) <= LineBuffer0(646);
            LineBuffer0(648) <= LineBuffer0(647);
            LineBuffer0(649) <= LineBuffer0(648);    
            LineBuffer0(650) <= LineBuffer0(649);
            LineBuffer0(651) <= LineBuffer0(650);
            LineBuffer0(652) <= LineBuffer0(651);
            LineBuffer0(653) <= LineBuffer0(652);
            LineBuffer0(654) <= LineBuffer0(653);
            LineBuffer0(655) <= LineBuffer0(654);
            LineBuffer0(656) <= LineBuffer0(655);
            LineBuffer0(657) <= LineBuffer0(656);
            LineBuffer0(658) <= LineBuffer0(657);
            LineBuffer0(659) <= LineBuffer0(658);    
            LineBuffer0(660) <= LineBuffer0(659);
            LineBuffer0(661) <= LineBuffer0(660);
            LineBuffer0(662) <= LineBuffer0(661);
            LineBuffer0(663) <= LineBuffer0(662);
            LineBuffer0(664) <= LineBuffer0(663);
            LineBuffer0(665) <= LineBuffer0(664);
            LineBuffer0(666) <= LineBuffer0(665);
            LineBuffer0(667) <= LineBuffer0(666);
            LineBuffer0(668) <= LineBuffer0(667);
            LineBuffer0(669) <= LineBuffer0(668);    
            LineBuffer0(670) <= LineBuffer0(669);
            LineBuffer0(671) <= LineBuffer0(670);
            LineBuffer0(672) <= LineBuffer0(671);
            LineBuffer0(673) <= LineBuffer0(672);
            LineBuffer0(674) <= LineBuffer0(673);
            LineBuffer0(675) <= LineBuffer0(674);
            LineBuffer0(676) <= LineBuffer0(675);
            LineBuffer0(677) <= LineBuffer0(676);
            LineBuffer0(678) <= LineBuffer0(677);
            LineBuffer0(679) <= LineBuffer0(678);    
            LineBuffer0(680) <= LineBuffer0(679);
            LineBuffer0(681) <= LineBuffer0(680);
            LineBuffer0(682) <= LineBuffer0(681);
            LineBuffer0(683) <= LineBuffer0(682);
            LineBuffer0(684) <= LineBuffer0(683);
            LineBuffer0(685) <= LineBuffer0(684);
            LineBuffer0(686) <= LineBuffer0(685);
            LineBuffer0(687) <= LineBuffer0(686);
            LineBuffer0(688) <= LineBuffer0(687);
            LineBuffer0(689) <= LineBuffer0(688);    
            LineBuffer0(690) <= LineBuffer0(689);
            LineBuffer0(691) <= LineBuffer0(690);
            LineBuffer0(692) <= LineBuffer0(691);
            LineBuffer0(693) <= LineBuffer0(692);
            LineBuffer0(694) <= LineBuffer0(693);
            LineBuffer0(695) <= LineBuffer0(694);
            LineBuffer0(696) <= LineBuffer0(695);
            LineBuffer0(697) <= LineBuffer0(696);
            LineBuffer0(698) <= LineBuffer0(697);
            LineBuffer0(699) <= LineBuffer0(698);    
            LineBuffer0(700) <= LineBuffer0(699);
            LineBuffer0(701) <= LineBuffer0(700);
            LineBuffer0(702) <= LineBuffer0(701);
            LineBuffer0(703) <= LineBuffer0(702);
            LineBuffer0(704) <= LineBuffer0(703);
            LineBuffer0(705) <= LineBuffer0(704);
            LineBuffer0(706) <= LineBuffer0(705);
            LineBuffer0(707) <= LineBuffer0(706);
            LineBuffer0(708) <= LineBuffer0(707);
            LineBuffer0(709) <= LineBuffer0(708);    
            LineBuffer0(710) <= LineBuffer0(709);
            LineBuffer0(711) <= LineBuffer0(710);
            LineBuffer0(712) <= LineBuffer0(711);
            LineBuffer0(713) <= LineBuffer0(712);
            LineBuffer0(714) <= LineBuffer0(713);
            LineBuffer0(715) <= LineBuffer0(714);
            LineBuffer0(716) <= LineBuffer0(715);
            LineBuffer0(717) <= LineBuffer0(716);
            LineBuffer0(718) <= LineBuffer0(717);
            LineBuffer0(719) <= LineBuffer0(718);    
            LineBuffer0(720) <= LineBuffer0(719);
            LineBuffer0(721) <= LineBuffer0(720);
            LineBuffer0(722) <= LineBuffer0(721);
            LineBuffer0(723) <= LineBuffer0(722);
            LineBuffer0(724) <= LineBuffer0(723);
            LineBuffer0(725) <= LineBuffer0(724);
            LineBuffer0(726) <= LineBuffer0(725);
            LineBuffer0(727) <= LineBuffer0(726);
            LineBuffer0(728) <= LineBuffer0(727);
            LineBuffer0(729) <= LineBuffer0(728);    
            LineBuffer0(730) <= LineBuffer0(729);
            LineBuffer0(731) <= LineBuffer0(730);
            LineBuffer0(732) <= LineBuffer0(731);
            LineBuffer0(733) <= LineBuffer0(732);
            LineBuffer0(734) <= LineBuffer0(733);
            LineBuffer0(735) <= LineBuffer0(734);
            LineBuffer0(736) <= LineBuffer0(735);
            LineBuffer0(737) <= LineBuffer0(736);
            LineBuffer0(738) <= LineBuffer0(737);
            LineBuffer0(739) <= LineBuffer0(738);    
            LineBuffer0(740) <= LineBuffer0(739);
            LineBuffer0(741) <= LineBuffer0(740);
            LineBuffer0(742) <= LineBuffer0(741);
            LineBuffer0(743) <= LineBuffer0(742);
            LineBuffer0(744) <= LineBuffer0(743);
            LineBuffer0(745) <= LineBuffer0(744);
            LineBuffer0(746) <= LineBuffer0(745);
            LineBuffer0(747) <= LineBuffer0(746);
            LineBuffer0(748) <= LineBuffer0(747);
            LineBuffer0(749) <= LineBuffer0(748);    
            LineBuffer0(750) <= LineBuffer0(749);
            LineBuffer0(751) <= LineBuffer0(750);
            LineBuffer0(752) <= LineBuffer0(751);
            LineBuffer0(753) <= LineBuffer0(752);
            LineBuffer0(754) <= LineBuffer0(753);
            LineBuffer0(755) <= LineBuffer0(754);
            LineBuffer0(756) <= LineBuffer0(755);
            LineBuffer0(757) <= LineBuffer0(756);
            LineBuffer0(758) <= LineBuffer0(757);
            LineBuffer0(759) <= LineBuffer0(758);    
            LineBuffer0(760) <= LineBuffer0(759);
            LineBuffer0(761) <= LineBuffer0(760);
            LineBuffer0(762) <= LineBuffer0(761);
            LineBuffer0(763) <= LineBuffer0(762);
            LineBuffer0(764) <= LineBuffer0(763);
            LineBuffer0(765) <= LineBuffer0(764);
            LineBuffer0(766) <= LineBuffer0(765);
            LineBuffer0(767) <= LineBuffer0(766);
            LineBuffer0(768) <= LineBuffer0(767);
            LineBuffer0(769) <= LineBuffer0(768);    
            LineBuffer0(770) <= LineBuffer0(769);
            LineBuffer0(771) <= LineBuffer0(770);
            LineBuffer0(772) <= LineBuffer0(771);
            LineBuffer0(773) <= LineBuffer0(772);
            LineBuffer0(774) <= LineBuffer0(773);
            LineBuffer0(775) <= LineBuffer0(774);
            LineBuffer0(776) <= LineBuffer0(775);
            LineBuffer0(777) <= LineBuffer0(776);
            LineBuffer0(778) <= LineBuffer0(777);
            LineBuffer0(779) <= LineBuffer0(778);    
            LineBuffer0(780) <= LineBuffer0(779);
            LineBuffer0(781) <= LineBuffer0(780);
            LineBuffer0(782) <= LineBuffer0(781);
            LineBuffer0(783) <= LineBuffer0(782);
            LineBuffer0(784) <= LineBuffer0(783);
            LineBuffer0(785) <= LineBuffer0(784);
            LineBuffer0(786) <= LineBuffer0(785);
            LineBuffer0(787) <= LineBuffer0(786);
            LineBuffer0(788) <= LineBuffer0(787);
            LineBuffer0(789) <= LineBuffer0(788);    
            LineBuffer0(790) <= LineBuffer0(789);
            LineBuffer0(791) <= LineBuffer0(790);
            LineBuffer0(792) <= LineBuffer0(791);
            LineBuffer0(793) <= LineBuffer0(792);
            LineBuffer0(794) <= LineBuffer0(793);
            LineBuffer0(795) <= LineBuffer0(794);
            LineBuffer0(796) <= LineBuffer0(795);
            LineBuffer0(797) <= LineBuffer0(796);
            LineBuffer0(798) <= LineBuffer0(797);
            LineBuffer0(799) <= LineBuffer0(798);    
            LineBuffer0(800) <= LineBuffer0(799);
            LineBuffer0(801) <= LineBuffer0(800);
            LineBuffer0(802) <= LineBuffer0(801);
            LineBuffer0(803) <= LineBuffer0(802);
            LineBuffer0(804) <= LineBuffer0(803);
            LineBuffer0(805) <= LineBuffer0(804);
            LineBuffer0(806) <= LineBuffer0(805);
            LineBuffer0(807) <= LineBuffer0(806);
            LineBuffer0(808) <= LineBuffer0(807);
            LineBuffer0(809) <= LineBuffer0(808);    
            LineBuffer0(810) <= LineBuffer0(809);
            LineBuffer0(811) <= LineBuffer0(810);
            LineBuffer0(812) <= LineBuffer0(811);
            LineBuffer0(813) <= LineBuffer0(812);
            LineBuffer0(814) <= LineBuffer0(813);
            LineBuffer0(815) <= LineBuffer0(814);
            LineBuffer0(816) <= LineBuffer0(815);
            LineBuffer0(817) <= LineBuffer0(816);
            LineBuffer0(818) <= LineBuffer0(817);
            LineBuffer0(819) <= LineBuffer0(818);    
            LineBuffer0(820) <= LineBuffer0(819);
            LineBuffer0(821) <= LineBuffer0(820);
            LineBuffer0(822) <= LineBuffer0(821);
            LineBuffer0(823) <= LineBuffer0(822);
            LineBuffer0(824) <= LineBuffer0(823);
            LineBuffer0(825) <= LineBuffer0(824);
            LineBuffer0(826) <= LineBuffer0(825);
            LineBuffer0(827) <= LineBuffer0(826);
            LineBuffer0(828) <= LineBuffer0(827);
            LineBuffer0(829) <= LineBuffer0(828);    
            LineBuffer0(830) <= LineBuffer0(829);
            LineBuffer0(831) <= LineBuffer0(830);
            LineBuffer0(832) <= LineBuffer0(831);
            LineBuffer0(833) <= LineBuffer0(832);
            LineBuffer0(834) <= LineBuffer0(833);
            LineBuffer0(835) <= LineBuffer0(834);
            LineBuffer0(836) <= LineBuffer0(835);
            LineBuffer0(837) <= LineBuffer0(836);
            LineBuffer0(838) <= LineBuffer0(837);
            LineBuffer0(839) <= LineBuffer0(838);
            LineBuffer0(840) <= LineBuffer0(839);
            LineBuffer0(841) <= LineBuffer0(840);
            LineBuffer0(842) <= LineBuffer0(841);
            LineBuffer0(843) <= LineBuffer0(842);
            LineBuffer0(844) <= LineBuffer0(843);
            LineBuffer0(845) <= LineBuffer0(844);
            LineBuffer0(846) <= LineBuffer0(845);
            LineBuffer0(847) <= LineBuffer0(846);
            LineBuffer0(848) <= LineBuffer0(847);
            LineBuffer0(849) <= LineBuffer0(848);    
            LineBuffer0(850) <= LineBuffer0(849);
            LineBuffer0(851) <= LineBuffer0(850);
            LineBuffer0(852) <= LineBuffer0(851);
            LineBuffer0(853) <= LineBuffer0(852);
            LineBuffer0(854) <= LineBuffer0(853);
            LineBuffer0(855) <= LineBuffer0(854);
            LineBuffer0(856) <= LineBuffer0(855);
            LineBuffer0(857) <= LineBuffer0(856);
            LineBuffer0(858) <= LineBuffer0(857);
            LineBuffer0(859) <= LineBuffer0(858);    
            LineBuffer0(860) <= LineBuffer0(859);
            LineBuffer0(861) <= LineBuffer0(860);
            LineBuffer0(862) <= LineBuffer0(861);
            LineBuffer0(863) <= LineBuffer0(862);
            LineBuffer0(864) <= LineBuffer0(863);
            LineBuffer0(865) <= LineBuffer0(864);
            LineBuffer0(866) <= LineBuffer0(865);
            LineBuffer0(867) <= LineBuffer0(866);
            LineBuffer0(868) <= LineBuffer0(867);
            LineBuffer0(869) <= LineBuffer0(868);    
            LineBuffer0(870) <= LineBuffer0(869);
            LineBuffer0(871) <= LineBuffer0(870);
            LineBuffer0(872) <= LineBuffer0(871);
            LineBuffer0(873) <= LineBuffer0(872);
            LineBuffer0(874) <= LineBuffer0(873);
            LineBuffer0(875) <= LineBuffer0(874);
            LineBuffer0(876) <= LineBuffer0(875);
            LineBuffer0(877) <= LineBuffer0(876);
            LineBuffer0(878) <= LineBuffer0(877);
            LineBuffer0(879) <= LineBuffer0(878);    
            LineBuffer0(880) <= LineBuffer0(879);
            LineBuffer0(881) <= LineBuffer0(880);
            LineBuffer0(882) <= LineBuffer0(881);
            LineBuffer0(883) <= LineBuffer0(882);
            LineBuffer0(884) <= LineBuffer0(883);
            LineBuffer0(885) <= LineBuffer0(884);
            LineBuffer0(886) <= LineBuffer0(885);
            LineBuffer0(887) <= LineBuffer0(886);
            LineBuffer0(888) <= LineBuffer0(887);
            LineBuffer0(889) <= LineBuffer0(888);    
            LineBuffer0(890) <= LineBuffer0(889);
            LineBuffer0(891) <= LineBuffer0(890);
            LineBuffer0(892) <= LineBuffer0(891);
            LineBuffer0(893) <= LineBuffer0(892);
            LineBuffer0(894) <= LineBuffer0(893);
            LineBuffer0(895) <= LineBuffer0(894);
            LineBuffer0(896) <= LineBuffer0(895);
            LineBuffer0(897) <= LineBuffer0(896);
            LineBuffer0(898) <= LineBuffer0(897);
            LineBuffer0(899) <= LineBuffer0(898);    
            LineBuffer0(900) <= LineBuffer0(899);
            LineBuffer0(901) <= LineBuffer0(900);
            LineBuffer0(902) <= LineBuffer0(901);
            LineBuffer0(903) <= LineBuffer0(902);
            LineBuffer0(904) <= LineBuffer0(903);
            LineBuffer0(905) <= LineBuffer0(904);
            LineBuffer0(906) <= LineBuffer0(905);
            LineBuffer0(907) <= LineBuffer0(906);
            LineBuffer0(908) <= LineBuffer0(907);
            LineBuffer0(909) <= LineBuffer0(908);    
            LineBuffer0(910) <= LineBuffer0(909);
            LineBuffer0(911) <= LineBuffer0(910);
            LineBuffer0(912) <= LineBuffer0(911);
            LineBuffer0(913) <= LineBuffer0(912);
            LineBuffer0(914) <= LineBuffer0(913);
            LineBuffer0(915) <= LineBuffer0(914);
            LineBuffer0(916) <= LineBuffer0(915);
            LineBuffer0(917) <= LineBuffer0(916);
            LineBuffer0(918) <= LineBuffer0(917);
            LineBuffer0(919) <= LineBuffer0(918);    
            LineBuffer0(920) <= LineBuffer0(919);
            LineBuffer0(921) <= LineBuffer0(920);
            LineBuffer0(922) <= LineBuffer0(921);
            LineBuffer0(923) <= LineBuffer0(922);
            LineBuffer0(924) <= LineBuffer0(923);
            LineBuffer0(925) <= LineBuffer0(924);
            LineBuffer0(926) <= LineBuffer0(925);
            LineBuffer0(927) <= LineBuffer0(926);
            LineBuffer0(928) <= LineBuffer0(927);
            LineBuffer0(929) <= LineBuffer0(928);    
            LineBuffer0(930) <= LineBuffer0(929);
            LineBuffer0(931) <= LineBuffer0(930);
            LineBuffer0(932) <= LineBuffer0(931);
            LineBuffer0(933) <= LineBuffer0(932);
            LineBuffer0(934) <= LineBuffer0(933);
            LineBuffer0(935) <= LineBuffer0(934);
            LineBuffer0(936) <= LineBuffer0(935);
            LineBuffer0(937) <= LineBuffer0(936);
            LineBuffer0(938) <= LineBuffer0(937);
            LineBuffer0(939) <= LineBuffer0(938);
            LineBuffer0(940) <= LineBuffer0(939);
            LineBuffer0(941) <= LineBuffer0(940);
            LineBuffer0(942) <= LineBuffer0(941);
            LineBuffer0(943) <= LineBuffer0(942);
            LineBuffer0(944) <= LineBuffer0(943);
            LineBuffer0(945) <= LineBuffer0(944);
            LineBuffer0(946) <= LineBuffer0(945);
            LineBuffer0(947) <= LineBuffer0(946);
            LineBuffer0(948) <= LineBuffer0(947);
            LineBuffer0(949) <= LineBuffer0(948);    
            LineBuffer0(950) <= LineBuffer0(949);
            LineBuffer0(951) <= LineBuffer0(950);
            LineBuffer0(952) <= LineBuffer0(951);
            LineBuffer0(953) <= LineBuffer0(952);
            LineBuffer0(954) <= LineBuffer0(953);
            LineBuffer0(955) <= LineBuffer0(954);
            LineBuffer0(956) <= LineBuffer0(955);
            LineBuffer0(957) <= LineBuffer0(956);
            LineBuffer0(958) <= LineBuffer0(957);
            LineBuffer0(959) <= LineBuffer0(958);    
            LineBuffer0(960) <= LineBuffer0(959);
            LineBuffer0(961) <= LineBuffer0(960);
            LineBuffer0(962) <= LineBuffer0(961);
            LineBuffer0(963) <= LineBuffer0(962);
            LineBuffer0(964) <= LineBuffer0(963);
            LineBuffer0(965) <= LineBuffer0(964);
            LineBuffer0(966) <= LineBuffer0(965);
            LineBuffer0(967) <= LineBuffer0(966);
            LineBuffer0(968) <= LineBuffer0(967);
            LineBuffer0(969) <= LineBuffer0(968);    
            LineBuffer0(970) <= LineBuffer0(969);
            LineBuffer0(971) <= LineBuffer0(970);
            LineBuffer0(972) <= LineBuffer0(971);
            LineBuffer0(973) <= LineBuffer0(972);
            LineBuffer0(974) <= LineBuffer0(973);
            LineBuffer0(975) <= LineBuffer0(974);
            LineBuffer0(976) <= LineBuffer0(975);
            LineBuffer0(977) <= LineBuffer0(976);
            LineBuffer0(978) <= LineBuffer0(977);
            LineBuffer0(979) <= LineBuffer0(978);    
            LineBuffer0(980) <= LineBuffer0(979);
            LineBuffer0(981) <= LineBuffer0(980);
            LineBuffer0(982) <= LineBuffer0(981);
            LineBuffer0(983) <= LineBuffer0(982);
            LineBuffer0(984) <= LineBuffer0(983);
            LineBuffer0(985) <= LineBuffer0(984);
            LineBuffer0(986) <= LineBuffer0(985);
            LineBuffer0(987) <= LineBuffer0(986);
            LineBuffer0(988) <= LineBuffer0(987);
            LineBuffer0(989) <= LineBuffer0(988);    
            LineBuffer0(990) <= LineBuffer0(989);
            LineBuffer0(991) <= LineBuffer0(990);
            LineBuffer0(992) <= LineBuffer0(991);
            LineBuffer0(993) <= LineBuffer0(992);
            LineBuffer0(994) <= LineBuffer0(993);
            LineBuffer0(995) <= LineBuffer0(994);
            LineBuffer0(996) <= LineBuffer0(995);
            LineBuffer0(997) <= LineBuffer0(996);
            LineBuffer0(998) <= LineBuffer0(997);
            LineBuffer0(999) <= LineBuffer0(998);    
            LineBuffer0(1000) <= LineBuffer0(999);
            LineBuffer0(1001) <= LineBuffer0(1000);
            LineBuffer0(1002) <= LineBuffer0(1001);
            LineBuffer0(1003) <= LineBuffer0(1002);
            LineBuffer0(1004) <= LineBuffer0(1003);
            LineBuffer0(1005) <= LineBuffer0(1004);
            LineBuffer0(1006) <= LineBuffer0(1005);
            LineBuffer0(1007) <= LineBuffer0(1006);
            LineBuffer0(1008) <= LineBuffer0(1007);
            LineBuffer0(1009) <= LineBuffer0(1008);    
            LineBuffer0(1010) <= LineBuffer0(1009);
            LineBuffer0(1011) <= LineBuffer0(1010);
            LineBuffer0(1012) <= LineBuffer0(1011);
            LineBuffer0(1013) <= LineBuffer0(1012);
            LineBuffer0(1014) <= LineBuffer0(1013);
            LineBuffer0(1015) <= LineBuffer0(1014);
            LineBuffer0(1016) <= LineBuffer0(1015);
            LineBuffer0(1017) <= LineBuffer0(1016);
            LineBuffer0(1018) <= LineBuffer0(1017);
            LineBuffer0(1019) <= LineBuffer0(1018);    
            LineBuffer0(1020) <= LineBuffer0(1019);
            LineBuffer0(1021) <= LineBuffer0(1020);
            LineBuffer0(1022) <= LineBuffer0(1021);
            LineBuffer0(1023) <= LineBuffer0(1022);
            LineBuffer0(1024) <= LineBuffer0(1023);
            LineBuffer0(1025) <= LineBuffer0(1024);
            LineBuffer0(1026) <= LineBuffer0(1025);
            LineBuffer0(1027) <= LineBuffer0(1026);
            LineBuffer0(1028) <= LineBuffer0(1027);
            LineBuffer0(1029) <= LineBuffer0(1028);    
            LineBuffer0(1030) <= LineBuffer0(1029);
            LineBuffer0(1031) <= LineBuffer0(1030);
            LineBuffer0(1032) <= LineBuffer0(1031);
            LineBuffer0(1033) <= LineBuffer0(1032);
            LineBuffer0(1034) <= LineBuffer0(1033);
            LineBuffer0(1035) <= LineBuffer0(1034);
            LineBuffer0(1036) <= LineBuffer0(1035);
            LineBuffer0(1037) <= LineBuffer0(1036);
            LineBuffer0(1038) <= LineBuffer0(1037);
            LineBuffer0(1039) <= LineBuffer0(1038);
            LineBuffer0(1040) <= LineBuffer0(1039);
            LineBuffer0(1041) <= LineBuffer0(1040);
            LineBuffer0(1042) <= LineBuffer0(1041);
            LineBuffer0(1043) <= LineBuffer0(1042);
            LineBuffer0(1044) <= LineBuffer0(1043);
            LineBuffer0(1045) <= LineBuffer0(1044);
            LineBuffer0(1046) <= LineBuffer0(1045);
            LineBuffer0(1047) <= LineBuffer0(1046);
            LineBuffer0(1048) <= LineBuffer0(1047);
            LineBuffer0(1049) <= LineBuffer0(1048);    
            LineBuffer0(1050) <= LineBuffer0(1049);
            LineBuffer0(1051) <= LineBuffer0(1050);
            LineBuffer0(1052) <= LineBuffer0(1051);
            LineBuffer0(1053) <= LineBuffer0(1052);
            LineBuffer0(1054) <= LineBuffer0(1053);
            LineBuffer0(1055) <= LineBuffer0(1054);
            LineBuffer0(1056) <= LineBuffer0(1055);
            LineBuffer0(1057) <= LineBuffer0(1056);
            LineBuffer0(1058) <= LineBuffer0(1057);
            LineBuffer0(1059) <= LineBuffer0(1058);    
            LineBuffer0(1060) <= LineBuffer0(1059);
            LineBuffer0(1061) <= LineBuffer0(1060);
            LineBuffer0(1062) <= LineBuffer0(1061);
            LineBuffer0(1063) <= LineBuffer0(1062);
            LineBuffer0(1064) <= LineBuffer0(1063);
            LineBuffer0(1065) <= LineBuffer0(1064);
            LineBuffer0(1066) <= LineBuffer0(1065);
            LineBuffer0(1067) <= LineBuffer0(1066);
            LineBuffer0(1068) <= LineBuffer0(1067);
            LineBuffer0(1069) <= LineBuffer0(1068);    
            LineBuffer0(1070) <= LineBuffer0(1069);
            LineBuffer0(1071) <= LineBuffer0(1070);
            LineBuffer0(1072) <= LineBuffer0(1071);
            LineBuffer0(1073) <= LineBuffer0(1072);
            LineBuffer0(1074) <= LineBuffer0(1073);
            LineBuffer0(1075) <= LineBuffer0(1074);
            LineBuffer0(1076) <= LineBuffer0(1075);
            LineBuffer0(1077) <= LineBuffer0(1076);
            LineBuffer0(1078) <= LineBuffer0(1077);
            LineBuffer0(1079) <= LineBuffer0(1078);    
            LineBuffer0(1080) <= LineBuffer0(1079);
            LineBuffer0(1081) <= LineBuffer0(1080);
            LineBuffer0(1082) <= LineBuffer0(1081);
            LineBuffer0(1083) <= LineBuffer0(1082);
            LineBuffer0(1084) <= LineBuffer0(1083);
            LineBuffer0(1085) <= LineBuffer0(1084);
            LineBuffer0(1086) <= LineBuffer0(1085);
            LineBuffer0(1087) <= LineBuffer0(1086);
            LineBuffer0(1088) <= LineBuffer0(1087);
            LineBuffer0(1089) <= LineBuffer0(1088);    
            LineBuffer0(1090) <= LineBuffer0(1089);
            LineBuffer0(1091) <= LineBuffer0(1090);
            LineBuffer0(1092) <= LineBuffer0(1091);
            LineBuffer0(1093) <= LineBuffer0(1092);
            LineBuffer0(1094) <= LineBuffer0(1093);
            LineBuffer0(1095) <= LineBuffer0(1094);
            LineBuffer0(1096) <= LineBuffer0(1095);
            LineBuffer0(1097) <= LineBuffer0(1096);
            LineBuffer0(1098) <= LineBuffer0(1097);
            LineBuffer0(1099) <= LineBuffer0(1098);    
            LineBuffer0(1100) <= LineBuffer0(1099);
            LineBuffer0(1101) <= LineBuffer0(1100);
            LineBuffer0(1102) <= LineBuffer0(1101);
            LineBuffer0(1103) <= LineBuffer0(1102);
            LineBuffer0(1104) <= LineBuffer0(1103);
            LineBuffer0(1105) <= LineBuffer0(1104);
            LineBuffer0(1106) <= LineBuffer0(1105);
            LineBuffer0(1107) <= LineBuffer0(1106);
            LineBuffer0(1108) <= LineBuffer0(1107);
            LineBuffer0(1109) <= LineBuffer0(1108);    
            LineBuffer0(1110) <= LineBuffer0(1109);
            LineBuffer0(1111) <= LineBuffer0(1110);
            LineBuffer0(1112) <= LineBuffer0(1111);
            LineBuffer0(1113) <= LineBuffer0(1112);
            LineBuffer0(1114) <= LineBuffer0(1113);
            LineBuffer0(1115) <= LineBuffer0(1114);
            LineBuffer0(1116) <= LineBuffer0(1115);
            LineBuffer0(1117) <= LineBuffer0(1116);
            LineBuffer0(1118) <= LineBuffer0(1117);
            LineBuffer0(1119) <= LineBuffer0(1118);    
            LineBuffer0(1120) <= LineBuffer0(1119);
            LineBuffer0(1121) <= LineBuffer0(1120);
            LineBuffer0(1122) <= LineBuffer0(1121);
            LineBuffer0(1123) <= LineBuffer0(1122);
            LineBuffer0(1124) <= LineBuffer0(1123);
            LineBuffer0(1125) <= LineBuffer0(1124);
            LineBuffer0(1126) <= LineBuffer0(1125);
            LineBuffer0(1127) <= LineBuffer0(1126);
            LineBuffer0(1128) <= LineBuffer0(1127);
            LineBuffer0(1129) <= LineBuffer0(1128);    
            LineBuffer0(1130) <= LineBuffer0(1129);
            LineBuffer0(1131) <= LineBuffer0(1130);
            LineBuffer0(1132) <= LineBuffer0(1131);
            LineBuffer0(1133) <= LineBuffer0(1132);
            LineBuffer0(1134) <= LineBuffer0(1133);
            LineBuffer0(1135) <= LineBuffer0(1134);
            LineBuffer0(1136) <= LineBuffer0(1135);
            LineBuffer0(1137) <= LineBuffer0(1136);
            LineBuffer0(1138) <= LineBuffer0(1137);
            LineBuffer0(1139) <= LineBuffer0(1138);
            LineBuffer0(1140) <= LineBuffer0(1139);
            LineBuffer0(1141) <= LineBuffer0(1140);
            LineBuffer0(1142) <= LineBuffer0(1141);
            LineBuffer0(1143) <= LineBuffer0(1142);
            LineBuffer0(1144) <= LineBuffer0(1143);
            LineBuffer0(1145) <= LineBuffer0(1144);
            LineBuffer0(1146) <= LineBuffer0(1145);
            LineBuffer0(1147) <= LineBuffer0(1146);
            LineBuffer0(1148) <= LineBuffer0(1147);
            LineBuffer0(1149) <= LineBuffer0(1148);    
            LineBuffer0(1150) <= LineBuffer0(1149);
            LineBuffer0(1151) <= LineBuffer0(1150);
            LineBuffer0(1152) <= LineBuffer0(1151);
            LineBuffer0(1153) <= LineBuffer0(1152);
            LineBuffer0(1154) <= LineBuffer0(1153);
            LineBuffer0(1155) <= LineBuffer0(1154);
            LineBuffer0(1156) <= LineBuffer0(1155);
            LineBuffer0(1157) <= LineBuffer0(1156);
            LineBuffer0(1158) <= LineBuffer0(1157);
            LineBuffer0(1159) <= LineBuffer0(1158);    
            LineBuffer0(1160) <= LineBuffer0(1159);
            LineBuffer0(1161) <= LineBuffer0(1160);
            LineBuffer0(1162) <= LineBuffer0(1161);
            LineBuffer0(1163) <= LineBuffer0(1162);
            LineBuffer0(1164) <= LineBuffer0(1163);
            LineBuffer0(1165) <= LineBuffer0(1164);
            LineBuffer0(1166) <= LineBuffer0(1165);
            LineBuffer0(1167) <= LineBuffer0(1166);
            LineBuffer0(1168) <= LineBuffer0(1167);
            LineBuffer0(1169) <= LineBuffer0(1168);    
            LineBuffer0(1170) <= LineBuffer0(1169);
            LineBuffer0(1171) <= LineBuffer0(1170);
            LineBuffer0(1172) <= LineBuffer0(1171);
            LineBuffer0(1173) <= LineBuffer0(1172);
            LineBuffer0(1174) <= LineBuffer0(1173);
            LineBuffer0(1175) <= LineBuffer0(1174);
            LineBuffer0(1176) <= LineBuffer0(1175);
            LineBuffer0(1177) <= LineBuffer0(1176);
            LineBuffer0(1178) <= LineBuffer0(1177);
            LineBuffer0(1179) <= LineBuffer0(1178);    
            LineBuffer0(1180) <= LineBuffer0(1179);
            LineBuffer0(1181) <= LineBuffer0(1180);
            LineBuffer0(1182) <= LineBuffer0(1181);
            LineBuffer0(1183) <= LineBuffer0(1182);
            LineBuffer0(1184) <= LineBuffer0(1183);
            LineBuffer0(1185) <= LineBuffer0(1184);
            LineBuffer0(1186) <= LineBuffer0(1185);
            LineBuffer0(1187) <= LineBuffer0(1186);
            LineBuffer0(1188) <= LineBuffer0(1187);
            LineBuffer0(1189) <= LineBuffer0(1188);    
            LineBuffer0(1190) <= LineBuffer0(1189);
            LineBuffer0(1191) <= LineBuffer0(1190);
            LineBuffer0(1192) <= LineBuffer0(1191);
            LineBuffer0(1193) <= LineBuffer0(1192);
            LineBuffer0(1194) <= LineBuffer0(1193);
            LineBuffer0(1195) <= LineBuffer0(1194);
            LineBuffer0(1196) <= LineBuffer0(1195);
            LineBuffer0(1197) <= LineBuffer0(1196);
            LineBuffer0(1198) <= LineBuffer0(1197);
            LineBuffer0(1199) <= LineBuffer0(1198);    
            LineBuffer0(1200) <= LineBuffer0(1199);
            LineBuffer0(1201) <= LineBuffer0(1200);
            LineBuffer0(1202) <= LineBuffer0(1201);
            LineBuffer0(1203) <= LineBuffer0(1202);
            LineBuffer0(1204) <= LineBuffer0(1203);
            LineBuffer0(1205) <= LineBuffer0(1204);
            LineBuffer0(1206) <= LineBuffer0(1205);
            LineBuffer0(1207) <= LineBuffer0(1206);
            LineBuffer0(1208) <= LineBuffer0(1207);
            LineBuffer0(1209) <= LineBuffer0(1208);    
            LineBuffer0(1210) <= LineBuffer0(1209);
            LineBuffer0(1211) <= LineBuffer0(1210);
            LineBuffer0(1212) <= LineBuffer0(1211);
            LineBuffer0(1213) <= LineBuffer0(1212);
            LineBuffer0(1214) <= LineBuffer0(1213);
            LineBuffer0(1215) <= LineBuffer0(1214);
            LineBuffer0(1216) <= LineBuffer0(1215);
            LineBuffer0(1217) <= LineBuffer0(1216);
            LineBuffer0(1218) <= LineBuffer0(1217);
            LineBuffer0(1219) <= LineBuffer0(1218);    
            LineBuffer0(1220) <= LineBuffer0(1219);
            LineBuffer0(1221) <= LineBuffer0(1220);
            LineBuffer0(1222) <= LineBuffer0(1221);
            LineBuffer0(1223) <= LineBuffer0(1222);
            LineBuffer0(1224) <= LineBuffer0(1223);
            LineBuffer0(1225) <= LineBuffer0(1224);
            LineBuffer0(1226) <= LineBuffer0(1225);
            LineBuffer0(1227) <= LineBuffer0(1226);
            LineBuffer0(1228) <= LineBuffer0(1227);
            LineBuffer0(1229) <= LineBuffer0(1228);    
            LineBuffer0(1230) <= LineBuffer0(1229);
            LineBuffer0(1231) <= LineBuffer0(1230);
            LineBuffer0(1232) <= LineBuffer0(1231);
            LineBuffer0(1233) <= LineBuffer0(1232);
            LineBuffer0(1234) <= LineBuffer0(1233);
            LineBuffer0(1235) <= LineBuffer0(1234);
            LineBuffer0(1236) <= LineBuffer0(1235);
            LineBuffer0(1237) <= LineBuffer0(1236);
            LineBuffer0(1238) <= LineBuffer0(1237);
            LineBuffer0(1239) <= LineBuffer0(1238);
            LineBuffer0(1240) <= LineBuffer0(1239);
            LineBuffer0(1241) <= LineBuffer0(1240);
            LineBuffer0(1242) <= LineBuffer0(1241);
            LineBuffer0(1243) <= LineBuffer0(1242);
            LineBuffer0(1244) <= LineBuffer0(1243);
            LineBuffer0(1245) <= LineBuffer0(1244);
            LineBuffer0(1246) <= LineBuffer0(1245);
            LineBuffer0(1247) <= LineBuffer0(1246);
            LineBuffer0(1248) <= LineBuffer0(1247);
            LineBuffer0(1249) <= LineBuffer0(1248);    
            LineBuffer0(1250) <= LineBuffer0(1249);
            LineBuffer0(1251) <= LineBuffer0(1250);
            LineBuffer0(1252) <= LineBuffer0(1251);
            LineBuffer0(1253) <= LineBuffer0(1252);
            LineBuffer0(1254) <= LineBuffer0(1253);
            LineBuffer0(1255) <= LineBuffer0(1254);
            LineBuffer0(1256) <= LineBuffer0(1255);
            LineBuffer0(1257) <= LineBuffer0(1256);
            LineBuffer0(1258) <= LineBuffer0(1257);
            LineBuffer0(1259) <= LineBuffer0(1258);    
            LineBuffer0(1260) <= LineBuffer0(1259);
            LineBuffer0(1261) <= LineBuffer0(1260);
            LineBuffer0(1262) <= LineBuffer0(1261);
            LineBuffer0(1263) <= LineBuffer0(1262);
            LineBuffer0(1264) <= LineBuffer0(1263);
            LineBuffer0(1265) <= LineBuffer0(1264);
            LineBuffer0(1266) <= LineBuffer0(1265);
            LineBuffer0(1267) <= LineBuffer0(1266);
            LineBuffer0(1268) <= LineBuffer0(1267);
            LineBuffer0(1269) <= LineBuffer0(1268);    
            LineBuffer0(1270) <= LineBuffer0(1269);
            LineBuffer0(1271) <= LineBuffer0(1270);
            LineBuffer0(1272) <= LineBuffer0(1271);
            LineBuffer0(1273) <= LineBuffer0(1272);
            LineBuffer0(1274) <= LineBuffer0(1273);
            LineBuffer0(1275) <= LineBuffer0(1274);
            LineBuffer0(1276) <= LineBuffer0(1275);
            LineBuffer0(1277) <= LineBuffer0(1276);
            LineBuffer0(1278) <= LineBuffer0(1277);
            LineBuffer0(1279) <= LineBuffer0(1278);
--            LineBuffer0(1280) <= LineBuffer0(1279);
--            LineBuffer0(1281) <= LineBuffer0(1280);
--            LineBuffer0(1282) <= LineBuffer0(1281);
--            LineBuffer0(1283) <= LineBuffer0(1282);
--            LineBuffer0(1284) <= LineBuffer0(1283);
--            LineBuffer0(1285) <= LineBuffer0(1284);
--            LineBuffer0(1286) <= LineBuffer0(1285);
--            LineBuffer0(1287) <= LineBuffer0(1286);
--            LineBuffer0(1288) <= LineBuffer0(1287);
--            LineBuffer0(1289) <= LineBuffer0(1288);    
--            LineBuffer0(1290) <= LineBuffer0(1289);
--            LineBuffer0(1291) <= LineBuffer0(1290);
--            LineBuffer0(1292) <= LineBuffer0(1291);
--            LineBuffer0(1293) <= LineBuffer0(1292);
--            LineBuffer0(1294) <= LineBuffer0(1293);
--            LineBuffer0(1295) <= LineBuffer0(1294);
--            LineBuffer0(1296) <= LineBuffer0(1295);
--            LineBuffer0(1297) <= LineBuffer0(1296);
--            LineBuffer0(1298) <= LineBuffer0(1297);
--            LineBuffer0(1299) <= LineBuffer0(1298);    
--            LineBuffer0(1300) <= LineBuffer0(1299);
--            LineBuffer0(1301) <= LineBuffer0(1300);
--            LineBuffer0(1302) <= LineBuffer0(1301);
--            LineBuffer0(1303) <= LineBuffer0(1302);
--            LineBuffer0(1304) <= LineBuffer0(1303);
--            LineBuffer0(1305) <= LineBuffer0(1304);
--            LineBuffer0(1306) <= LineBuffer0(1305);
--            LineBuffer0(1307) <= LineBuffer0(1306);
--            LineBuffer0(1308) <= LineBuffer0(1307);
--            LineBuffer0(1309) <= LineBuffer0(1308);    
--            LineBuffer0(1310) <= LineBuffer0(1309);
--            LineBuffer0(1311) <= LineBuffer0(1310);
--            LineBuffer0(1312) <= LineBuffer0(1311);
--            LineBuffer0(1313) <= LineBuffer0(1312);
--            LineBuffer0(1314) <= LineBuffer0(1313);
--            LineBuffer0(1315) <= LineBuffer0(1314);
--            LineBuffer0(1316) <= LineBuffer0(1315);
--            LineBuffer0(1317) <= LineBuffer0(1316);
--            LineBuffer0(1318) <= LineBuffer0(1317);
--            LineBuffer0(1319) <= LineBuffer0(1318);    
--            LineBuffer0(1320) <= LineBuffer0(1319);
--            LineBuffer0(1321) <= LineBuffer0(1320);
--            LineBuffer0(1322) <= LineBuffer0(1321);
--            LineBuffer0(1323) <= LineBuffer0(1322);
--            LineBuffer0(1324) <= LineBuffer0(1323);
--            LineBuffer0(1325) <= LineBuffer0(1324);
--            LineBuffer0(1326) <= LineBuffer0(1325);
--            LineBuffer0(1327) <= LineBuffer0(1326);
--            LineBuffer0(1328) <= LineBuffer0(1327);
--            LineBuffer0(1329) <= LineBuffer0(1328);    
--            LineBuffer0(1330) <= LineBuffer0(1329);
--            LineBuffer0(1331) <= LineBuffer0(1330);
--            LineBuffer0(1332) <= LineBuffer0(1331);
--            LineBuffer0(1333) <= LineBuffer0(1332);
--            LineBuffer0(1334) <= LineBuffer0(1333);
--            LineBuffer0(1335) <= LineBuffer0(1334);
--            LineBuffer0(1336) <= LineBuffer0(1335);
--            LineBuffer0(1337) <= LineBuffer0(1336);
--            LineBuffer0(1338) <= LineBuffer0(1337);
--            LineBuffer0(1339) <= LineBuffer0(1338);    
--            LineBuffer0(1340) <= LineBuffer0(1339);
--            LineBuffer0(1341) <= LineBuffer0(1340);
--            LineBuffer0(1342) <= LineBuffer0(1341);
--            LineBuffer0(1343) <= LineBuffer0(1342);
--            LineBuffer0(1344) <= LineBuffer0(1343);
--            LineBuffer0(1345) <= LineBuffer0(1344);
--            LineBuffer0(1346) <= LineBuffer0(1345);
--            LineBuffer0(1347) <= LineBuffer0(1346);
--            LineBuffer0(1348) <= LineBuffer0(1347);
--            LineBuffer0(1349) <= LineBuffer0(1348);    
--            LineBuffer0(1350) <= LineBuffer0(1349);
--            LineBuffer0(1351) <= LineBuffer0(1350);
--            LineBuffer0(1352) <= LineBuffer0(1351);
--            LineBuffer0(1353) <= LineBuffer0(1352);
--            LineBuffer0(1354) <= LineBuffer0(1353);
--            LineBuffer0(1355) <= LineBuffer0(1354);
--            LineBuffer0(1356) <= LineBuffer0(1355);
--            LineBuffer0(1357) <= LineBuffer0(1356);
--            LineBuffer0(1358) <= LineBuffer0(1357);
--            LineBuffer0(1359) <= LineBuffer0(1358);    
--            LineBuffer0(1360) <= LineBuffer0(1359);
--            LineBuffer0(1361) <= LineBuffer0(1360);
--            LineBuffer0(1362) <= LineBuffer0(1361);
--            LineBuffer0(1363) <= LineBuffer0(1362);
--            LineBuffer0(1364) <= LineBuffer0(1363);
--            LineBuffer0(1365) <= LineBuffer0(1364);
--            LineBuffer0(1366) <= LineBuffer0(1365);
--            LineBuffer0(1367) <= LineBuffer0(1366);
--            LineBuffer0(1368) <= LineBuffer0(1367);
--            LineBuffer0(1369) <= LineBuffer0(1368);    
--            LineBuffer0(1370) <= LineBuffer0(1369);
--            LineBuffer0(1371) <= LineBuffer0(1370);
--            LineBuffer0(1372) <= LineBuffer0(1371);
--            LineBuffer0(1373) <= LineBuffer0(1372);
--            LineBuffer0(1374) <= LineBuffer0(1373);
--            LineBuffer0(1375) <= LineBuffer0(1374);
--            LineBuffer0(1376) <= LineBuffer0(1375);
--            LineBuffer0(1377) <= LineBuffer0(1376);
--            LineBuffer0(1378) <= LineBuffer0(1377);
--            LineBuffer0(1379) <= LineBuffer0(1378);    
--            LineBuffer0(1380) <= LineBuffer0(1379);
--            LineBuffer0(1381) <= LineBuffer0(1380);
--            LineBuffer0(1382) <= LineBuffer0(1381);
--            LineBuffer0(1383) <= LineBuffer0(1382);
--            LineBuffer0(1384) <= LineBuffer0(1383);
--            LineBuffer0(1385) <= LineBuffer0(1384);
--            LineBuffer0(1386) <= LineBuffer0(1385);
--            LineBuffer0(1387) <= LineBuffer0(1386);
--            LineBuffer0(1388) <= LineBuffer0(1387);
--            LineBuffer0(1389) <= LineBuffer0(1388);    
--            LineBuffer0(1390) <= LineBuffer0(1389);
--            LineBuffer0(1391) <= LineBuffer0(1390);
--            LineBuffer0(1392) <= LineBuffer0(1391);
--            LineBuffer0(1393) <= LineBuffer0(1392);
--            LineBuffer0(1394) <= LineBuffer0(1393);
--            LineBuffer0(1395) <= LineBuffer0(1394);
--            LineBuffer0(1396) <= LineBuffer0(1395);
--            LineBuffer0(1397) <= LineBuffer0(1396);
--            LineBuffer0(1398) <= LineBuffer0(1397);
--            LineBuffer0(1399) <= LineBuffer0(1398);    
--            LineBuffer0(1400) <= LineBuffer0(1399);
--            LineBuffer0(1401) <= LineBuffer0(1400);
--            LineBuffer0(1402) <= LineBuffer0(1401);
--            LineBuffer0(1403) <= LineBuffer0(1402);
--            LineBuffer0(1404) <= LineBuffer0(1403);
--            LineBuffer0(1405) <= LineBuffer0(1404);
--            LineBuffer0(1406) <= LineBuffer0(1405);
--            LineBuffer0(1407) <= LineBuffer0(1406);
--            LineBuffer0(1408) <= LineBuffer0(1407);
--            LineBuffer0(1409) <= LineBuffer0(1408);    
--            LineBuffer0(1410) <= LineBuffer0(1409);
--            LineBuffer0(1411) <= LineBuffer0(1410);
--            LineBuffer0(1412) <= LineBuffer0(1411);
--            LineBuffer0(1413) <= LineBuffer0(1412);
--            LineBuffer0(1414) <= LineBuffer0(1413);
--            LineBuffer0(1415) <= LineBuffer0(1414);
--            LineBuffer0(1416) <= LineBuffer0(1415);
--            LineBuffer0(1417) <= LineBuffer0(1416);
--            LineBuffer0(1418) <= LineBuffer0(1417);
--            LineBuffer0(1419) <= LineBuffer0(1418);    
--            LineBuffer0(1420) <= LineBuffer0(1419);
--            LineBuffer0(1421) <= LineBuffer0(1420);
--            LineBuffer0(1422) <= LineBuffer0(1421);
--            LineBuffer0(1423) <= LineBuffer0(1422);
--            LineBuffer0(1424) <= LineBuffer0(1423);
--            LineBuffer0(1425) <= LineBuffer0(1424);
--            LineBuffer0(1426) <= LineBuffer0(1425);
--            LineBuffer0(1427) <= LineBuffer0(1426);
--            LineBuffer0(1428) <= LineBuffer0(1427);
--            LineBuffer0(1429) <= LineBuffer0(1428);    
--            LineBuffer0(1430) <= LineBuffer0(1429);
--            LineBuffer0(1431) <= LineBuffer0(1430);
--            LineBuffer0(1432) <= LineBuffer0(1431);
--            LineBuffer0(1433) <= LineBuffer0(1432);
--            LineBuffer0(1434) <= LineBuffer0(1433);
--            LineBuffer0(1435) <= LineBuffer0(1434);
--            LineBuffer0(1436) <= LineBuffer0(1435);
--            LineBuffer0(1437) <= LineBuffer0(1436);
--            LineBuffer0(1438) <= LineBuffer0(1437);
--            LineBuffer0(1439) <= LineBuffer0(1438);    
--            LineBuffer0(1440) <= LineBuffer0(1439);
--            LineBuffer0(1441) <= LineBuffer0(1440);
--            LineBuffer0(1442) <= LineBuffer0(1441);
--            LineBuffer0(1443) <= LineBuffer0(1442);
--            LineBuffer0(1444) <= LineBuffer0(1443);
--            LineBuffer0(1445) <= LineBuffer0(1444);
--            LineBuffer0(1446) <= LineBuffer0(1445);
--            LineBuffer0(1447) <= LineBuffer0(1446);
--            LineBuffer0(1448) <= LineBuffer0(1447);
--            LineBuffer0(1449) <= LineBuffer0(1448);    
--            LineBuffer0(1450) <= LineBuffer0(1449);
--            LineBuffer0(1451) <= LineBuffer0(1450);
--            LineBuffer0(1452) <= LineBuffer0(1451);
--            LineBuffer0(1453) <= LineBuffer0(1452);
--            LineBuffer0(1454) <= LineBuffer0(1453);
--            LineBuffer0(1455) <= LineBuffer0(1454);
--            LineBuffer0(1456) <= LineBuffer0(1455);
--            LineBuffer0(1457) <= LineBuffer0(1456);
--            LineBuffer0(1458) <= LineBuffer0(1457);
--            LineBuffer0(1459) <= LineBuffer0(1458);    
--            LineBuffer0(1460) <= LineBuffer0(1459);
--            LineBuffer0(1461) <= LineBuffer0(1460);
--            LineBuffer0(1462) <= LineBuffer0(1461);
--            LineBuffer0(1463) <= LineBuffer0(1462);
--            LineBuffer0(1464) <= LineBuffer0(1463);
--            LineBuffer0(1465) <= LineBuffer0(1464);
--            LineBuffer0(1466) <= LineBuffer0(1465);
--            LineBuffer0(1467) <= LineBuffer0(1466);
--            LineBuffer0(1468) <= LineBuffer0(1467);
--            LineBuffer0(1469) <= LineBuffer0(1468);    
--            LineBuffer0(1470) <= LineBuffer0(1469);
--            LineBuffer0(1471) <= LineBuffer0(1470);
--            LineBuffer0(1472) <= LineBuffer0(1471);
--            LineBuffer0(1473) <= LineBuffer0(1472);
--            LineBuffer0(1474) <= LineBuffer0(1473);
--            LineBuffer0(1475) <= LineBuffer0(1474);
--            LineBuffer0(1476) <= LineBuffer0(1475);
--            LineBuffer0(1477) <= LineBuffer0(1476);
--            LineBuffer0(1478) <= LineBuffer0(1477);
--            LineBuffer0(1479) <= LineBuffer0(1478);
--            LineBuffer0(1480) <= LineBuffer0(1479);
--            LineBuffer0(1481) <= LineBuffer0(1480);
--            LineBuffer0(1482) <= LineBuffer0(1481);
--            LineBuffer0(1483) <= LineBuffer0(1482);
--            LineBuffer0(1484) <= LineBuffer0(1483);
--            LineBuffer0(1485) <= LineBuffer0(1484);
--            LineBuffer0(1486) <= LineBuffer0(1485);
--            LineBuffer0(1487) <= LineBuffer0(1486);
--            LineBuffer0(1488) <= LineBuffer0(1487);
--            LineBuffer0(1489) <= LineBuffer0(1488);    
--            LineBuffer0(1490) <= LineBuffer0(1489);
--            LineBuffer0(1491) <= LineBuffer0(1490);
--            LineBuffer0(1492) <= LineBuffer0(1491);
--            LineBuffer0(1493) <= LineBuffer0(1492);
--            LineBuffer0(1494) <= LineBuffer0(1493);
--            LineBuffer0(1495) <= LineBuffer0(1494);
--            LineBuffer0(1496) <= LineBuffer0(1495);
--            LineBuffer0(1497) <= LineBuffer0(1496);
--            LineBuffer0(1498) <= LineBuffer0(1497);
--            LineBuffer0(1499) <= LineBuffer0(1498);    
--            LineBuffer0(1500) <= LineBuffer0(1499);
--            LineBuffer0(1501) <= LineBuffer0(1500);
--            LineBuffer0(1502) <= LineBuffer0(1501);
--            LineBuffer0(1503) <= LineBuffer0(1502);
--            LineBuffer0(1504) <= LineBuffer0(1503);
--            LineBuffer0(1505) <= LineBuffer0(1504);
--            LineBuffer0(1506) <= LineBuffer0(1505);
--            LineBuffer0(1507) <= LineBuffer0(1506);
--            LineBuffer0(1508) <= LineBuffer0(1507);
--            LineBuffer0(1509) <= LineBuffer0(1508);    
--            LineBuffer0(1510) <= LineBuffer0(1509);
--            LineBuffer0(1511) <= LineBuffer0(1510);
--            LineBuffer0(1512) <= LineBuffer0(1511);
--            LineBuffer0(1513) <= LineBuffer0(1512);
--            LineBuffer0(1514) <= LineBuffer0(1513);
--            LineBuffer0(1515) <= LineBuffer0(1514);
--            LineBuffer0(1516) <= LineBuffer0(1515);
--            LineBuffer0(1517) <= LineBuffer0(1516);
--            LineBuffer0(1518) <= LineBuffer0(1517);
--            LineBuffer0(1519) <= LineBuffer0(1518);    
--            LineBuffer0(1520) <= LineBuffer0(1519);
--            LineBuffer0(1521) <= LineBuffer0(1520);
--            LineBuffer0(1522) <= LineBuffer0(1521);
--            LineBuffer0(1523) <= LineBuffer0(1522);
--            LineBuffer0(1524) <= LineBuffer0(1523);
--            LineBuffer0(1525) <= LineBuffer0(1524);
--            LineBuffer0(1526) <= LineBuffer0(1525);
--            LineBuffer0(1527) <= LineBuffer0(1526);
--            LineBuffer0(1528) <= LineBuffer0(1527);
--            LineBuffer0(1529) <= LineBuffer0(1528);    
--            LineBuffer0(1530) <= LineBuffer0(1529);
--            LineBuffer0(1531) <= LineBuffer0(1530);
--            LineBuffer0(1532) <= LineBuffer0(1531);
--            LineBuffer0(1533) <= LineBuffer0(1532);
--            LineBuffer0(1534) <= LineBuffer0(1533);
--            LineBuffer0(1535) <= LineBuffer0(1534);
--            LineBuffer0(1536) <= LineBuffer0(1535);
--            LineBuffer0(1537) <= LineBuffer0(1536);
--            LineBuffer0(1538) <= LineBuffer0(1537);
--            LineBuffer0(1539) <= LineBuffer0(1538);    
--            LineBuffer0(1540) <= LineBuffer0(1539);
--            LineBuffer0(1541) <= LineBuffer0(1540);
--            LineBuffer0(1542) <= LineBuffer0(1541);
--            LineBuffer0(1543) <= LineBuffer0(1542);
--            LineBuffer0(1544) <= LineBuffer0(1543);
--            LineBuffer0(1545) <= LineBuffer0(1544);
--            LineBuffer0(1546) <= LineBuffer0(1545);
--            LineBuffer0(1547) <= LineBuffer0(1546);
--            LineBuffer0(1548) <= LineBuffer0(1547);
--            LineBuffer0(1549) <= LineBuffer0(1548);    
--            LineBuffer0(1550) <= LineBuffer0(1549);
--            LineBuffer0(1551) <= LineBuffer0(1550);
--            LineBuffer0(1552) <= LineBuffer0(1551);
--            LineBuffer0(1553) <= LineBuffer0(1552);
--            LineBuffer0(1554) <= LineBuffer0(1553);
--            LineBuffer0(1555) <= LineBuffer0(1554);
--            LineBuffer0(1556) <= LineBuffer0(1555);
--            LineBuffer0(1557) <= LineBuffer0(1556);
--            LineBuffer0(1558) <= LineBuffer0(1557);
--            LineBuffer0(1559) <= LineBuffer0(1558);    
--            LineBuffer0(1560) <= LineBuffer0(1559);
--            LineBuffer0(1561) <= LineBuffer0(1560);
--            LineBuffer0(1562) <= LineBuffer0(1561);
--            LineBuffer0(1563) <= LineBuffer0(1562);
--            LineBuffer0(1564) <= LineBuffer0(1563);
--            LineBuffer0(1565) <= LineBuffer0(1564);
--            LineBuffer0(1566) <= LineBuffer0(1565);
--            LineBuffer0(1567) <= LineBuffer0(1566);
--            LineBuffer0(1568) <= LineBuffer0(1567);
--            LineBuffer0(1569) <= LineBuffer0(1568);    
--            LineBuffer0(1570) <= LineBuffer0(1569);
--            LineBuffer0(1571) <= LineBuffer0(1570);
--            LineBuffer0(1572) <= LineBuffer0(1571);
--            LineBuffer0(1573) <= LineBuffer0(1572);
--            LineBuffer0(1574) <= LineBuffer0(1573);
--            LineBuffer0(1575) <= LineBuffer0(1574);
--            LineBuffer0(1576) <= LineBuffer0(1575);
--            LineBuffer0(1577) <= LineBuffer0(1576);
--            LineBuffer0(1578) <= LineBuffer0(1577);
--            LineBuffer0(1579) <= LineBuffer0(1578);
--            LineBuffer0(1580) <= LineBuffer0(1579);
--            LineBuffer0(1581) <= LineBuffer0(1580);
--            LineBuffer0(1582) <= LineBuffer0(1581);
--            LineBuffer0(1583) <= LineBuffer0(1582);
--            LineBuffer0(1584) <= LineBuffer0(1583);
--            LineBuffer0(1585) <= LineBuffer0(1584);
--            LineBuffer0(1586) <= LineBuffer0(1585);
--            LineBuffer0(1587) <= LineBuffer0(1586);
--            LineBuffer0(1588) <= LineBuffer0(1587);
--            LineBuffer0(1589) <= LineBuffer0(1588);    
--            LineBuffer0(1590) <= LineBuffer0(1589);
--            LineBuffer0(1591) <= LineBuffer0(1590);
--            LineBuffer0(1592) <= LineBuffer0(1591);
--            LineBuffer0(1593) <= LineBuffer0(1592);
--            LineBuffer0(1594) <= LineBuffer0(1593);
--            LineBuffer0(1595) <= LineBuffer0(1594);
--            LineBuffer0(1596) <= LineBuffer0(1595);
--            LineBuffer0(1597) <= LineBuffer0(1596);
--            LineBuffer0(1598) <= LineBuffer0(1597);
--            LineBuffer0(1599) <= LineBuffer0(1598);    
--            LineBuffer0(1600) <= LineBuffer0(1599);
--            LineBuffer0(1601) <= LineBuffer0(1600);
--            LineBuffer0(1602) <= LineBuffer0(1601);
--            LineBuffer0(1603) <= LineBuffer0(1602);
--            LineBuffer0(1604) <= LineBuffer0(1603);
--            LineBuffer0(1605) <= LineBuffer0(1604);
--            LineBuffer0(1606) <= LineBuffer0(1605);
--            LineBuffer0(1607) <= LineBuffer0(1606);
--            LineBuffer0(1608) <= LineBuffer0(1607);
--            LineBuffer0(1609) <= LineBuffer0(1608);    
--            LineBuffer0(1610) <= LineBuffer0(1609);
--            LineBuffer0(1611) <= LineBuffer0(1610);
--            LineBuffer0(1612) <= LineBuffer0(1611);
--            LineBuffer0(1613) <= LineBuffer0(1612);
--            LineBuffer0(1614) <= LineBuffer0(1613);
--            LineBuffer0(1615) <= LineBuffer0(1614);
--            LineBuffer0(1616) <= LineBuffer0(1615);
--            LineBuffer0(1617) <= LineBuffer0(1616);
--            LineBuffer0(1618) <= LineBuffer0(1617);
--            LineBuffer0(1619) <= LineBuffer0(1618);    
--            LineBuffer0(1620) <= LineBuffer0(1619);
--            LineBuffer0(1621) <= LineBuffer0(1620);
--            LineBuffer0(1622) <= LineBuffer0(1621);
--            LineBuffer0(1623) <= LineBuffer0(1622);
--            LineBuffer0(1624) <= LineBuffer0(1623);
--            LineBuffer0(1625) <= LineBuffer0(1624);
--            LineBuffer0(1626) <= LineBuffer0(1625);
--            LineBuffer0(1627) <= LineBuffer0(1626);
--            LineBuffer0(1628) <= LineBuffer0(1627);
--            LineBuffer0(1629) <= LineBuffer0(1628);    
--            LineBuffer0(1630) <= LineBuffer0(1629);
--            LineBuffer0(1631) <= LineBuffer0(1630);
--            LineBuffer0(1632) <= LineBuffer0(1631);
--            LineBuffer0(1633) <= LineBuffer0(1632);
--            LineBuffer0(1634) <= LineBuffer0(1633);
--            LineBuffer0(1635) <= LineBuffer0(1634);
--            LineBuffer0(1636) <= LineBuffer0(1635);
--            LineBuffer0(1637) <= LineBuffer0(1636);
--            LineBuffer0(1638) <= LineBuffer0(1637);
--            LineBuffer0(1639) <= LineBuffer0(1638);    
--            LineBuffer0(1640) <= LineBuffer0(1639);
--            LineBuffer0(1641) <= LineBuffer0(1640);
--            LineBuffer0(1642) <= LineBuffer0(1641);
--            LineBuffer0(1643) <= LineBuffer0(1642);
--            LineBuffer0(1644) <= LineBuffer0(1643);
--            LineBuffer0(1645) <= LineBuffer0(1644);
--            LineBuffer0(1646) <= LineBuffer0(1645);
--            LineBuffer0(1647) <= LineBuffer0(1646);
--            LineBuffer0(1648) <= LineBuffer0(1647);
--            LineBuffer0(1649) <= LineBuffer0(1648);    
--            LineBuffer0(1650) <= LineBuffer0(1649);
--            LineBuffer0(1651) <= LineBuffer0(1650);
--            LineBuffer0(1652) <= LineBuffer0(1651);
--            LineBuffer0(1653) <= LineBuffer0(1652);
--            LineBuffer0(1654) <= LineBuffer0(1653);
--            LineBuffer0(1655) <= LineBuffer0(1654);
--            LineBuffer0(1656) <= LineBuffer0(1655);
--            LineBuffer0(1657) <= LineBuffer0(1656);
--            LineBuffer0(1658) <= LineBuffer0(1657);
--            LineBuffer0(1659) <= LineBuffer0(1658);    
--            LineBuffer0(1660) <= LineBuffer0(1659);
--            LineBuffer0(1661) <= LineBuffer0(1660);
--            LineBuffer0(1662) <= LineBuffer0(1661);
--            LineBuffer0(1663) <= LineBuffer0(1662);
--            LineBuffer0(1664) <= LineBuffer0(1663);
--            LineBuffer0(1665) <= LineBuffer0(1664);
--            LineBuffer0(1666) <= LineBuffer0(1665);
--            LineBuffer0(1667) <= LineBuffer0(1666);
--            LineBuffer0(1668) <= LineBuffer0(1667);
--            LineBuffer0(1669) <= LineBuffer0(1668);    
--            LineBuffer0(1670) <= LineBuffer0(1669);
--            LineBuffer0(1671) <= LineBuffer0(1670);
--            LineBuffer0(1672) <= LineBuffer0(1671);
--            LineBuffer0(1673) <= LineBuffer0(1672);
--            LineBuffer0(1674) <= LineBuffer0(1673);
--            LineBuffer0(1675) <= LineBuffer0(1674);
--            LineBuffer0(1676) <= LineBuffer0(1675);
--            LineBuffer0(1677) <= LineBuffer0(1676);
--            LineBuffer0(1678) <= LineBuffer0(1677);
--            LineBuffer0(1679) <= LineBuffer0(1678);
--            LineBuffer0(1680) <= LineBuffer0(1679);
--            LineBuffer0(1681) <= LineBuffer0(1680);
--            LineBuffer0(1682) <= LineBuffer0(1681);
--            LineBuffer0(1683) <= LineBuffer0(1682);
--            LineBuffer0(1684) <= LineBuffer0(1683);
--            LineBuffer0(1685) <= LineBuffer0(1684);
--            LineBuffer0(1686) <= LineBuffer0(1685);
--            LineBuffer0(1687) <= LineBuffer0(1686);
--            LineBuffer0(1688) <= LineBuffer0(1687);
--            LineBuffer0(1689) <= LineBuffer0(1688);    
--            LineBuffer0(1690) <= LineBuffer0(1689);
--            LineBuffer0(1691) <= LineBuffer0(1690);
--            LineBuffer0(1692) <= LineBuffer0(1691);
--            LineBuffer0(1693) <= LineBuffer0(1692);
--            LineBuffer0(1694) <= LineBuffer0(1693);
--            LineBuffer0(1695) <= LineBuffer0(1694);
--            LineBuffer0(1696) <= LineBuffer0(1695);
--            LineBuffer0(1697) <= LineBuffer0(1696);
--            LineBuffer0(1698) <= LineBuffer0(1697);
--            LineBuffer0(1699) <= LineBuffer0(1698);    
--            LineBuffer0(1700) <= LineBuffer0(1699);
--            LineBuffer0(1701) <= LineBuffer0(1700);
--            LineBuffer0(1702) <= LineBuffer0(1701);
--            LineBuffer0(1703) <= LineBuffer0(1702);
--            LineBuffer0(1704) <= LineBuffer0(1703);
--            LineBuffer0(1705) <= LineBuffer0(1704);
--            LineBuffer0(1706) <= LineBuffer0(1705);
--            LineBuffer0(1707) <= LineBuffer0(1706);
--            LineBuffer0(1708) <= LineBuffer0(1707);
--            LineBuffer0(1709) <= LineBuffer0(1708);    
--            LineBuffer0(1710) <= LineBuffer0(1709);
--            LineBuffer0(1711) <= LineBuffer0(1710);
--            LineBuffer0(1712) <= LineBuffer0(1711);
--            LineBuffer0(1713) <= LineBuffer0(1712);
--            LineBuffer0(1714) <= LineBuffer0(1713);
--            LineBuffer0(1715) <= LineBuffer0(1714);
--            LineBuffer0(1716) <= LineBuffer0(1715);
--            LineBuffer0(1717) <= LineBuffer0(1716);
--            LineBuffer0(1718) <= LineBuffer0(1717);
--            LineBuffer0(1719) <= LineBuffer0(1718);    
--            LineBuffer0(1720) <= LineBuffer0(1719);
--            LineBuffer0(1721) <= LineBuffer0(1720);
--            LineBuffer0(1722) <= LineBuffer0(1721);
--            LineBuffer0(1723) <= LineBuffer0(1722);
--            LineBuffer0(1724) <= LineBuffer0(1723);
--            LineBuffer0(1725) <= LineBuffer0(1724);
--            LineBuffer0(1726) <= LineBuffer0(1725);
--            LineBuffer0(1727) <= LineBuffer0(1726);
--            LineBuffer0(1728) <= LineBuffer0(1727);
--            LineBuffer0(1729) <= LineBuffer0(1728);    
--            LineBuffer0(1730) <= LineBuffer0(1729);
--            LineBuffer0(1731) <= LineBuffer0(1730);
--            LineBuffer0(1732) <= LineBuffer0(1731);
--            LineBuffer0(1733) <= LineBuffer0(1732);
--            LineBuffer0(1734) <= LineBuffer0(1733);
--            LineBuffer0(1735) <= LineBuffer0(1734);
--            LineBuffer0(1736) <= LineBuffer0(1735);
--            LineBuffer0(1737) <= LineBuffer0(1736);
--            LineBuffer0(1738) <= LineBuffer0(1737);
--            LineBuffer0(1739) <= LineBuffer0(1738);    
--            LineBuffer0(1740) <= LineBuffer0(1739);
--            LineBuffer0(1741) <= LineBuffer0(1740);
--            LineBuffer0(1742) <= LineBuffer0(1741);
--            LineBuffer0(1743) <= LineBuffer0(1742);
--            LineBuffer0(1744) <= LineBuffer0(1743);
--            LineBuffer0(1745) <= LineBuffer0(1744);
--            LineBuffer0(1746) <= LineBuffer0(1745);
--            LineBuffer0(1747) <= LineBuffer0(1746);
--            LineBuffer0(1748) <= LineBuffer0(1747);
--            LineBuffer0(1749) <= LineBuffer0(1748);    
--            LineBuffer0(1750) <= LineBuffer0(1749);
--            LineBuffer0(1751) <= LineBuffer0(1750);
--            LineBuffer0(1752) <= LineBuffer0(1751);
--            LineBuffer0(1753) <= LineBuffer0(1752);
--            LineBuffer0(1754) <= LineBuffer0(1753);
--            LineBuffer0(1755) <= LineBuffer0(1754);
--            LineBuffer0(1756) <= LineBuffer0(1755);
--            LineBuffer0(1757) <= LineBuffer0(1756);
--            LineBuffer0(1758) <= LineBuffer0(1757);
--            LineBuffer0(1759) <= LineBuffer0(1758);    
--            LineBuffer0(1760) <= LineBuffer0(1759);
--            LineBuffer0(1761) <= LineBuffer0(1760);
--            LineBuffer0(1762) <= LineBuffer0(1761);
--            LineBuffer0(1763) <= LineBuffer0(1762);
--            LineBuffer0(1764) <= LineBuffer0(1763);
--            LineBuffer0(1765) <= LineBuffer0(1764);
--            LineBuffer0(1766) <= LineBuffer0(1765);
--            LineBuffer0(1767) <= LineBuffer0(1766);
--            LineBuffer0(1768) <= LineBuffer0(1767);
--            LineBuffer0(1769) <= LineBuffer0(1768);    
--            LineBuffer0(1770) <= LineBuffer0(1769);
--            LineBuffer0(1771) <= LineBuffer0(1770);
--            LineBuffer0(1772) <= LineBuffer0(1771);
--            LineBuffer0(1773) <= LineBuffer0(1772);
--            LineBuffer0(1774) <= LineBuffer0(1773);
--            LineBuffer0(1775) <= LineBuffer0(1774);
--            LineBuffer0(1776) <= LineBuffer0(1775);
--            LineBuffer0(1777) <= LineBuffer0(1776);
--            LineBuffer0(1778) <= LineBuffer0(1777);
--            LineBuffer0(1779) <= LineBuffer0(1778);
--            LineBuffer0(1780) <= LineBuffer0(1779);
--            LineBuffer0(1781) <= LineBuffer0(1780);
--            LineBuffer0(1782) <= LineBuffer0(1781);
--            LineBuffer0(1783) <= LineBuffer0(1782);
--            LineBuffer0(1784) <= LineBuffer0(1783);
--            LineBuffer0(1785) <= LineBuffer0(1784);
--            LineBuffer0(1786) <= LineBuffer0(1785);
--            LineBuffer0(1787) <= LineBuffer0(1786);
--            LineBuffer0(1788) <= LineBuffer0(1787);
--            LineBuffer0(1789) <= LineBuffer0(1788);    
--            LineBuffer0(1790) <= LineBuffer0(1789);
--            LineBuffer0(1791) <= LineBuffer0(1790);
--            LineBuffer0(1792) <= LineBuffer0(1791);
--            LineBuffer0(1793) <= LineBuffer0(1792);
--            LineBuffer0(1794) <= LineBuffer0(1793);
--            LineBuffer0(1795) <= LineBuffer0(1794);
--            LineBuffer0(1796) <= LineBuffer0(1795);
--            LineBuffer0(1797) <= LineBuffer0(1796);
--            LineBuffer0(1798) <= LineBuffer0(1797);
--            LineBuffer0(1799) <= LineBuffer0(1798);    
--            LineBuffer0(1800) <= LineBuffer0(1799);
--            LineBuffer0(1801) <= LineBuffer0(1800);
--            LineBuffer0(1802) <= LineBuffer0(1801);
--            LineBuffer0(1803) <= LineBuffer0(1802);
--            LineBuffer0(1804) <= LineBuffer0(1803);
--            LineBuffer0(1805) <= LineBuffer0(1804);
--            LineBuffer0(1806) <= LineBuffer0(1805);
--            LineBuffer0(1807) <= LineBuffer0(1806);
--            LineBuffer0(1808) <= LineBuffer0(1807);
--            LineBuffer0(1809) <= LineBuffer0(1808);    
--            LineBuffer0(1810) <= LineBuffer0(1809);
--            LineBuffer0(1811) <= LineBuffer0(1810);
--            LineBuffer0(1812) <= LineBuffer0(1811);
--            LineBuffer0(1813) <= LineBuffer0(1812);
--            LineBuffer0(1814) <= LineBuffer0(1813);
--            LineBuffer0(1815) <= LineBuffer0(1814);
--            LineBuffer0(1816) <= LineBuffer0(1815);
--            LineBuffer0(1817) <= LineBuffer0(1816);
--            LineBuffer0(1818) <= LineBuffer0(1817);
--            LineBuffer0(1819) <= LineBuffer0(1818);    
--            LineBuffer0(1820) <= LineBuffer0(1819);
--            LineBuffer0(1821) <= LineBuffer0(1820);
--            LineBuffer0(1822) <= LineBuffer0(1821);
--            LineBuffer0(1823) <= LineBuffer0(1822);
--            LineBuffer0(1824) <= LineBuffer0(1823);
--            LineBuffer0(1825) <= LineBuffer0(1824);
--            LineBuffer0(1826) <= LineBuffer0(1825);
--            LineBuffer0(1827) <= LineBuffer0(1826);
--            LineBuffer0(1828) <= LineBuffer0(1827);
--            LineBuffer0(1829) <= LineBuffer0(1828);    
--            LineBuffer0(1830) <= LineBuffer0(1829);
--            LineBuffer0(1831) <= LineBuffer0(1830);
--            LineBuffer0(1832) <= LineBuffer0(1831);
--            LineBuffer0(1833) <= LineBuffer0(1832);
--            LineBuffer0(1834) <= LineBuffer0(1833);
--            LineBuffer0(1835) <= LineBuffer0(1834);
--            LineBuffer0(1836) <= LineBuffer0(1835);
--            LineBuffer0(1837) <= LineBuffer0(1836);
--            LineBuffer0(1838) <= LineBuffer0(1837);
--            LineBuffer0(1839) <= LineBuffer0(1838);    
--            LineBuffer0(1840) <= LineBuffer0(1839);
--            LineBuffer0(1841) <= LineBuffer0(1840);
--            LineBuffer0(1842) <= LineBuffer0(1841);
--            LineBuffer0(1843) <= LineBuffer0(1842);
--            LineBuffer0(1844) <= LineBuffer0(1843);
--            LineBuffer0(1845) <= LineBuffer0(1844);
--            LineBuffer0(1846) <= LineBuffer0(1845);
--            LineBuffer0(1847) <= LineBuffer0(1846);
--            LineBuffer0(1848) <= LineBuffer0(1847);
--            LineBuffer0(1849) <= LineBuffer0(1848);    
--            LineBuffer0(1850) <= LineBuffer0(1849);
--            LineBuffer0(1851) <= LineBuffer0(1850);
--            LineBuffer0(1852) <= LineBuffer0(1851);
--            LineBuffer0(1853) <= LineBuffer0(1852);
--            LineBuffer0(1854) <= LineBuffer0(1853);
--            LineBuffer0(1855) <= LineBuffer0(1854);
--            LineBuffer0(1856) <= LineBuffer0(1855);
--            LineBuffer0(1857) <= LineBuffer0(1856);
--            LineBuffer0(1858) <= LineBuffer0(1857);
--            LineBuffer0(1859) <= LineBuffer0(1858);    
--            LineBuffer0(1860) <= LineBuffer0(1859);
--            LineBuffer0(1861) <= LineBuffer0(1860);
--            LineBuffer0(1862) <= LineBuffer0(1861);
--            LineBuffer0(1863) <= LineBuffer0(1862);
--            LineBuffer0(1864) <= LineBuffer0(1863);
--            LineBuffer0(1865) <= LineBuffer0(1864);
--            LineBuffer0(1866) <= LineBuffer0(1865);
--            LineBuffer0(1867) <= LineBuffer0(1866);
--            LineBuffer0(1868) <= LineBuffer0(1867);
--            LineBuffer0(1869) <= LineBuffer0(1868);    
--            LineBuffer0(1870) <= LineBuffer0(1869);
--            LineBuffer0(1871) <= LineBuffer0(1870);
--            LineBuffer0(1872) <= LineBuffer0(1871);
--            LineBuffer0(1873) <= LineBuffer0(1872);
--            LineBuffer0(1874) <= LineBuffer0(1873);
--            LineBuffer0(1875) <= LineBuffer0(1874);
--            LineBuffer0(1876) <= LineBuffer0(1875);
--            LineBuffer0(1877) <= LineBuffer0(1876);
--            LineBuffer0(1878) <= LineBuffer0(1877);
--            LineBuffer0(1879) <= LineBuffer0(1878);
--            LineBuffer0(1880) <= LineBuffer0(1879);
--            LineBuffer0(1881) <= LineBuffer0(1880);
--            LineBuffer0(1882) <= LineBuffer0(1881);
--            LineBuffer0(1883) <= LineBuffer0(1882);
--            LineBuffer0(1884) <= LineBuffer0(1883);
--            LineBuffer0(1885) <= LineBuffer0(1884);
--            LineBuffer0(1886) <= LineBuffer0(1885);
--            LineBuffer0(1887) <= LineBuffer0(1886);
--            LineBuffer0(1888) <= LineBuffer0(1887);
--            LineBuffer0(1889) <= LineBuffer0(1888);    
--            LineBuffer0(1890) <= LineBuffer0(1889);
--            LineBuffer0(1891) <= LineBuffer0(1890);
--            LineBuffer0(1892) <= LineBuffer0(1891);
--            LineBuffer0(1893) <= LineBuffer0(1892);
--            LineBuffer0(1894) <= LineBuffer0(1893);
--            LineBuffer0(1895) <= LineBuffer0(1894);
--            LineBuffer0(1896) <= LineBuffer0(1895);
--            LineBuffer0(1897) <= LineBuffer0(1896);
--            LineBuffer0(1898) <= LineBuffer0(1897);
--            LineBuffer0(1899) <= LineBuffer0(1898);    
--            LineBuffer0(1900) <= LineBuffer0(1899);
--            LineBuffer0(1901) <= LineBuffer0(1900);
--            LineBuffer0(1902) <= LineBuffer0(1901);
--            LineBuffer0(1903) <= LineBuffer0(1902);
--            LineBuffer0(1904) <= LineBuffer0(1903);
--            LineBuffer0(1905) <= LineBuffer0(1904);
--            LineBuffer0(1906) <= LineBuffer0(1905);
--            LineBuffer0(1907) <= LineBuffer0(1906);
--            LineBuffer0(1908) <= LineBuffer0(1907);
--            LineBuffer0(1909) <= LineBuffer0(1908);    
--            LineBuffer0(1910) <= LineBuffer0(1909);
--            LineBuffer0(1911) <= LineBuffer0(1910);
--            LineBuffer0(1912) <= LineBuffer0(1911);
--            LineBuffer0(1913) <= LineBuffer0(1912);
--            LineBuffer0(1914) <= LineBuffer0(1913);
--            LineBuffer0(1915) <= LineBuffer0(1914);
--            LineBuffer0(1916) <= LineBuffer0(1915);
--            LineBuffer0(1917) <= LineBuffer0(1916);
--            LineBuffer0(1918) <= LineBuffer0(1917);
--            LineBuffer0(1919) <= LineBuffer0(1918);
		
		
			

			LineBuffer1(0) <= LineBuffer0(1279);
			LineBuffer1(1) <= LineBuffer1(0);
			LineBuffer1(2) <= LineBuffer1(1);
			LineBuffer1(3) <= LineBuffer1(2);
			LineBuffer1(4) <= LineBuffer1(3);
			LineBuffer1(5) <= LineBuffer1(4);
			LineBuffer1(6) <= LineBuffer1(5);
			LineBuffer1(7) <= LineBuffer1(6);
			LineBuffer1(8) <= LineBuffer1(7);
			LineBuffer1(9) <= LineBuffer1(8);	
			LineBuffer1(10) <= LineBuffer1(9);
			LineBuffer1(11) <= LineBuffer1(10);
			LineBuffer1(12) <= LineBuffer1(11);
			LineBuffer1(13) <= LineBuffer1(12);
			LineBuffer1(14) <= LineBuffer1(13);
			LineBuffer1(15) <= LineBuffer1(14);
			LineBuffer1(16) <= LineBuffer1(15);
			LineBuffer1(17) <= LineBuffer1(16);
			LineBuffer1(18) <= LineBuffer1(17);
			LineBuffer1(19) <= LineBuffer1(18);	
			LineBuffer1(20) <= LineBuffer1(19);
			LineBuffer1(21) <= LineBuffer1(20);
			LineBuffer1(22) <= LineBuffer1(21);
			LineBuffer1(23) <= LineBuffer1(22);
			LineBuffer1(24) <= LineBuffer1(23);
			LineBuffer1(25) <= LineBuffer1(24);
			LineBuffer1(26) <= LineBuffer1(25);
			LineBuffer1(27) <= LineBuffer1(26);
			LineBuffer1(28) <= LineBuffer1(27);
			LineBuffer1(29) <= LineBuffer1(28);	
			LineBuffer1(30) <= LineBuffer1(29);
			LineBuffer1(31) <= LineBuffer1(30);
			LineBuffer1(32) <= LineBuffer1(31);
			LineBuffer1(33) <= LineBuffer1(32);
			LineBuffer1(34) <= LineBuffer1(33);
			LineBuffer1(35) <= LineBuffer1(34);
			LineBuffer1(36) <= LineBuffer1(35);
			LineBuffer1(37) <= LineBuffer1(36);
			LineBuffer1(38) <= LineBuffer1(37);
			LineBuffer1(39) <= LineBuffer1(38);	
			LineBuffer1(40) <= LineBuffer1(39);
			LineBuffer1(41) <= LineBuffer1(40);
			LineBuffer1(42) <= LineBuffer1(41);
			LineBuffer1(43) <= LineBuffer1(42);
			LineBuffer1(44) <= LineBuffer1(43);
			LineBuffer1(45) <= LineBuffer1(44);
			LineBuffer1(46) <= LineBuffer1(45);
			LineBuffer1(47) <= LineBuffer1(46);
			LineBuffer1(48) <= LineBuffer1(47);
			LineBuffer1(49) <= LineBuffer1(48);	
			LineBuffer1(50) <= LineBuffer1(49);
			LineBuffer1(51) <= LineBuffer1(50);
			LineBuffer1(52) <= LineBuffer1(51);
			LineBuffer1(53) <= LineBuffer1(52);
			LineBuffer1(54) <= LineBuffer1(53);
			LineBuffer1(55) <= LineBuffer1(54);
			LineBuffer1(56) <= LineBuffer1(55);
			LineBuffer1(57) <= LineBuffer1(56);
			LineBuffer1(58) <= LineBuffer1(57);
			LineBuffer1(59) <= LineBuffer1(58);	
			LineBuffer1(60) <= LineBuffer1(59);
			LineBuffer1(61) <= LineBuffer1(60);
			LineBuffer1(62) <= LineBuffer1(61);
			LineBuffer1(63) <= LineBuffer1(62);
			LineBuffer1(64) <= LineBuffer1(63);
			LineBuffer1(65) <= LineBuffer1(64);
			LineBuffer1(66) <= LineBuffer1(65);
			LineBuffer1(67) <= LineBuffer1(66);
			LineBuffer1(68) <= LineBuffer1(67);
			LineBuffer1(69) <= LineBuffer1(68);	
			LineBuffer1(70) <= LineBuffer1(69);
			LineBuffer1(71) <= LineBuffer1(70);
			LineBuffer1(72) <= LineBuffer1(71);
			LineBuffer1(73) <= LineBuffer1(72);
			LineBuffer1(74) <= LineBuffer1(73);
			LineBuffer1(75) <= LineBuffer1(74);
			LineBuffer1(76) <= LineBuffer1(75);
			LineBuffer1(77) <= LineBuffer1(76);
			LineBuffer1(78) <= LineBuffer1(77);
			LineBuffer1(79) <= LineBuffer1(78);	
			LineBuffer1(80) <= LineBuffer1(79);
			LineBuffer1(81) <= LineBuffer1(80);
			LineBuffer1(82) <= LineBuffer1(81);
			LineBuffer1(83) <= LineBuffer1(82);
			LineBuffer1(84) <= LineBuffer1(83);
			LineBuffer1(85) <= LineBuffer1(84);
			LineBuffer1(86) <= LineBuffer1(85);
			LineBuffer1(87) <= LineBuffer1(86);
			LineBuffer1(88) <= LineBuffer1(87);
			LineBuffer1(89) <= LineBuffer1(88);	
			LineBuffer1(90) <= LineBuffer1(89);
			LineBuffer1(91) <= LineBuffer1(90);
			LineBuffer1(92) <= LineBuffer1(91);
			LineBuffer1(93) <= LineBuffer1(92);
			LineBuffer1(94) <= LineBuffer1(93);
			LineBuffer1(95) <= LineBuffer1(94);
			LineBuffer1(96) <= LineBuffer1(95);
			LineBuffer1(97) <= LineBuffer1(96);
			LineBuffer1(98) <= LineBuffer1(97);
			LineBuffer1(99) <= LineBuffer1(98);	
			LineBuffer1(100) <= LineBuffer1(99);
			LineBuffer1(101) <= LineBuffer1(100);
			LineBuffer1(102) <= LineBuffer1(101);
			LineBuffer1(103) <= LineBuffer1(102);
			LineBuffer1(104) <= LineBuffer1(103);
			LineBuffer1(105) <= LineBuffer1(104);
			LineBuffer1(106) <= LineBuffer1(105);
			LineBuffer1(107) <= LineBuffer1(106);
			LineBuffer1(108) <= LineBuffer1(107);
			LineBuffer1(109) <= LineBuffer1(108);	
			LineBuffer1(110) <= LineBuffer1(109);
			LineBuffer1(111) <= LineBuffer1(110);
			LineBuffer1(112) <= LineBuffer1(111);
			LineBuffer1(113) <= LineBuffer1(112);
			LineBuffer1(114) <= LineBuffer1(113);
			LineBuffer1(115) <= LineBuffer1(114);
			LineBuffer1(116) <= LineBuffer1(115);
			LineBuffer1(117) <= LineBuffer1(116);
			LineBuffer1(118) <= LineBuffer1(117);
			LineBuffer1(119) <= LineBuffer1(118);	
			LineBuffer1(120) <= LineBuffer1(119);
			LineBuffer1(121) <= LineBuffer1(120);
			LineBuffer1(122) <= LineBuffer1(121);
			LineBuffer1(123) <= LineBuffer1(122);
			LineBuffer1(124) <= LineBuffer1(123);
			LineBuffer1(125) <= LineBuffer1(124);
			LineBuffer1(126) <= LineBuffer1(125);
			LineBuffer1(127) <= LineBuffer1(126);
			LineBuffer1(128) <= LineBuffer1(127);
			LineBuffer1(129) <= LineBuffer1(128);	
			LineBuffer1(130) <= LineBuffer1(129);
			LineBuffer1(131) <= LineBuffer1(130);
			LineBuffer1(132) <= LineBuffer1(131);
			LineBuffer1(133) <= LineBuffer1(132);
			LineBuffer1(134) <= LineBuffer1(133);
			LineBuffer1(135) <= LineBuffer1(134);
			LineBuffer1(136) <= LineBuffer1(135);
			LineBuffer1(137) <= LineBuffer1(136);
			LineBuffer1(138) <= LineBuffer1(137);
			LineBuffer1(139) <= LineBuffer1(138);	
			LineBuffer1(140) <= LineBuffer1(139);
			LineBuffer1(141) <= LineBuffer1(140);
			LineBuffer1(142) <= LineBuffer1(141);
			LineBuffer1(143) <= LineBuffer1(142);
			LineBuffer1(144) <= LineBuffer1(143);
			LineBuffer1(145) <= LineBuffer1(144);
			LineBuffer1(146) <= LineBuffer1(145);
			LineBuffer1(147) <= LineBuffer1(146);
			LineBuffer1(148) <= LineBuffer1(147);
			LineBuffer1(149) <= LineBuffer1(148);	
			LineBuffer1(150) <= LineBuffer1(149);
			LineBuffer1(151) <= LineBuffer1(150);
			LineBuffer1(152) <= LineBuffer1(151);
			LineBuffer1(153) <= LineBuffer1(152);
			LineBuffer1(154) <= LineBuffer1(153);
			LineBuffer1(155) <= LineBuffer1(154);
			LineBuffer1(156) <= LineBuffer1(155);
			LineBuffer1(157) <= LineBuffer1(156);
			LineBuffer1(158) <= LineBuffer1(157);
			LineBuffer1(159) <= LineBuffer1(158);	
			LineBuffer1(160) <= LineBuffer1(159);
			LineBuffer1(161) <= LineBuffer1(160);
			LineBuffer1(162) <= LineBuffer1(161);
			LineBuffer1(163) <= LineBuffer1(162);
			LineBuffer1(164) <= LineBuffer1(163);
			LineBuffer1(165) <= LineBuffer1(164);
			LineBuffer1(166) <= LineBuffer1(165);
			LineBuffer1(167) <= LineBuffer1(166);
			LineBuffer1(168) <= LineBuffer1(167);
			LineBuffer1(169) <= LineBuffer1(168);	
			LineBuffer1(170) <= LineBuffer1(169);
			LineBuffer1(171) <= LineBuffer1(170);
			LineBuffer1(172) <= LineBuffer1(171);
			LineBuffer1(173) <= LineBuffer1(172);
			LineBuffer1(174) <= LineBuffer1(173);
			LineBuffer1(175) <= LineBuffer1(174);
			LineBuffer1(176) <= LineBuffer1(175);
			LineBuffer1(177) <= LineBuffer1(176);
			LineBuffer1(178) <= LineBuffer1(177);
			LineBuffer1(179) <= LineBuffer1(178);	
			LineBuffer1(180) <= LineBuffer1(179);
			LineBuffer1(181) <= LineBuffer1(180);
			LineBuffer1(182) <= LineBuffer1(181);
			LineBuffer1(183) <= LineBuffer1(182);
			LineBuffer1(184) <= LineBuffer1(183);
			LineBuffer1(185) <= LineBuffer1(184);
			LineBuffer1(186) <= LineBuffer1(185);
			LineBuffer1(187) <= LineBuffer1(186);
			LineBuffer1(188) <= LineBuffer1(187);
			LineBuffer1(189) <= LineBuffer1(188);	
			LineBuffer1(190) <= LineBuffer1(189);
			LineBuffer1(191) <= LineBuffer1(190);
			LineBuffer1(192) <= LineBuffer1(191);
			LineBuffer1(193) <= LineBuffer1(192);
			LineBuffer1(194) <= LineBuffer1(193);
			LineBuffer1(195) <= LineBuffer1(194);
			LineBuffer1(196) <= LineBuffer1(195);
			LineBuffer1(197) <= LineBuffer1(196);
			LineBuffer1(198) <= LineBuffer1(197);
			LineBuffer1(199) <= LineBuffer1(198);
			LineBuffer1(200) <= LineBuffer1(199);
			LineBuffer1(201) <= LineBuffer1(200);
			LineBuffer1(202) <= LineBuffer1(201);
			LineBuffer1(203) <= LineBuffer1(202);
			LineBuffer1(204) <= LineBuffer1(203);
			LineBuffer1(205) <= LineBuffer1(204);
			LineBuffer1(206) <= LineBuffer1(205);
			LineBuffer1(207) <= LineBuffer1(206);
			LineBuffer1(208) <= LineBuffer1(207);
			LineBuffer1(209) <= LineBuffer1(208);	
			LineBuffer1(210) <= LineBuffer1(209);
			LineBuffer1(211) <= LineBuffer1(210);
			LineBuffer1(212) <= LineBuffer1(211);
			LineBuffer1(213) <= LineBuffer1(212);
			LineBuffer1(214) <= LineBuffer1(213);
			LineBuffer1(215) <= LineBuffer1(214);
			LineBuffer1(216) <= LineBuffer1(215);
			LineBuffer1(217) <= LineBuffer1(216);
			LineBuffer1(218) <= LineBuffer1(217);
			LineBuffer1(219) <= LineBuffer1(218);	
			LineBuffer1(220) <= LineBuffer1(219);
			LineBuffer1(221) <= LineBuffer1(220);
			LineBuffer1(222) <= LineBuffer1(221);
			LineBuffer1(223) <= LineBuffer1(222);
			LineBuffer1(224) <= LineBuffer1(223);
			LineBuffer1(225) <= LineBuffer1(224);
			LineBuffer1(226) <= LineBuffer1(225);
			LineBuffer1(227) <= LineBuffer1(226);
			LineBuffer1(228) <= LineBuffer1(227);
			LineBuffer1(229) <= LineBuffer1(228);	
			LineBuffer1(230) <= LineBuffer1(229);
			LineBuffer1(231) <= LineBuffer1(230);
			LineBuffer1(232) <= LineBuffer1(231);
			LineBuffer1(233) <= LineBuffer1(232);
			LineBuffer1(234) <= LineBuffer1(233);
			LineBuffer1(235) <= LineBuffer1(234);
			LineBuffer1(236) <= LineBuffer1(235);
			LineBuffer1(237) <= LineBuffer1(236);
			LineBuffer1(238) <= LineBuffer1(237);
			LineBuffer1(239) <= LineBuffer1(238);	
			LineBuffer1(240) <= LineBuffer1(239);
			LineBuffer1(241) <= LineBuffer1(240);
			LineBuffer1(242) <= LineBuffer1(241);
			LineBuffer1(243) <= LineBuffer1(242);
			LineBuffer1(244) <= LineBuffer1(243);
			LineBuffer1(245) <= LineBuffer1(244);
			LineBuffer1(246) <= LineBuffer1(245);
			LineBuffer1(247) <= LineBuffer1(246);
			LineBuffer1(248) <= LineBuffer1(247);
			LineBuffer1(249) <= LineBuffer1(248);	
			LineBuffer1(250) <= LineBuffer1(249);
			LineBuffer1(251) <= LineBuffer1(250);
			LineBuffer1(252) <= LineBuffer1(251);
			LineBuffer1(253) <= LineBuffer1(252);
			LineBuffer1(254) <= LineBuffer1(253);
			LineBuffer1(255) <= LineBuffer1(254);
			LineBuffer1(256) <= LineBuffer1(255);
			LineBuffer1(257) <= LineBuffer1(256);
			LineBuffer1(258) <= LineBuffer1(257);
			LineBuffer1(259) <= LineBuffer1(258);	
			LineBuffer1(260) <= LineBuffer1(259);
			LineBuffer1(261) <= LineBuffer1(260);
			LineBuffer1(262) <= LineBuffer1(261);
			LineBuffer1(263) <= LineBuffer1(262);
			LineBuffer1(264) <= LineBuffer1(263);
			LineBuffer1(265) <= LineBuffer1(264);
			LineBuffer1(266) <= LineBuffer1(265);
			LineBuffer1(267) <= LineBuffer1(266);
			LineBuffer1(268) <= LineBuffer1(267);
			LineBuffer1(269) <= LineBuffer1(268);	
			LineBuffer1(270) <= LineBuffer1(269);
			LineBuffer1(271) <= LineBuffer1(270);
			LineBuffer1(272) <= LineBuffer1(271);
			LineBuffer1(273) <= LineBuffer1(272);
			LineBuffer1(274) <= LineBuffer1(273);
			LineBuffer1(275) <= LineBuffer1(274);
			LineBuffer1(276) <= LineBuffer1(275);
			LineBuffer1(277) <= LineBuffer1(276);
			LineBuffer1(278) <= LineBuffer1(277);
			LineBuffer1(279) <= LineBuffer1(278);	
			LineBuffer1(280) <= LineBuffer1(279);
			LineBuffer1(281) <= LineBuffer1(280);
			LineBuffer1(282) <= LineBuffer1(281);
			LineBuffer1(283) <= LineBuffer1(282);
			LineBuffer1(284) <= LineBuffer1(283);
			LineBuffer1(285) <= LineBuffer1(284);
			LineBuffer1(286) <= LineBuffer1(285);
			LineBuffer1(287) <= LineBuffer1(286);
			LineBuffer1(288) <= LineBuffer1(287);
			LineBuffer1(289) <= LineBuffer1(288);	
			LineBuffer1(290) <= LineBuffer1(289);
			LineBuffer1(291) <= LineBuffer1(290);
			LineBuffer1(292) <= LineBuffer1(291);
			LineBuffer1(293) <= LineBuffer1(292);
			LineBuffer1(294) <= LineBuffer1(293);
			LineBuffer1(295) <= LineBuffer1(294);
			LineBuffer1(296) <= LineBuffer1(295);
			LineBuffer1(297) <= LineBuffer1(296);
			LineBuffer1(298) <= LineBuffer1(297);
			LineBuffer1(299) <= LineBuffer1(298);	
			LineBuffer1(300) <= LineBuffer1(299);	
			LineBuffer1(301) <= LineBuffer1(300);
			LineBuffer1(302) <= LineBuffer1(301);
			LineBuffer1(303) <= LineBuffer1(302);
			LineBuffer1(304) <= LineBuffer1(303);
			LineBuffer1(305) <= LineBuffer1(304);
			LineBuffer1(306) <= LineBuffer1(305);
			LineBuffer1(307) <= LineBuffer1(306);
			LineBuffer1(308) <= LineBuffer1(307);
			LineBuffer1(309) <= LineBuffer1(308);	
			LineBuffer1(310) <= LineBuffer1(309);
			LineBuffer1(311) <= LineBuffer1(310);
			LineBuffer1(312) <= LineBuffer1(311);
			LineBuffer1(313) <= LineBuffer1(312);
			LineBuffer1(314) <= LineBuffer1(313);
			LineBuffer1(315) <= LineBuffer1(314);
			LineBuffer1(316) <= LineBuffer1(315);
			LineBuffer1(317) <= LineBuffer1(316);
			LineBuffer1(318) <= LineBuffer1(317);
			LineBuffer1(319) <= LineBuffer1(318);	
			LineBuffer1(320) <= LineBuffer1(319);
			LineBuffer1(321) <= LineBuffer1(320);
			LineBuffer1(322) <= LineBuffer1(321);
			LineBuffer1(323) <= LineBuffer1(322);
			LineBuffer1(324) <= LineBuffer1(323);
			LineBuffer1(325) <= LineBuffer1(324);
			LineBuffer1(326) <= LineBuffer1(325);
			LineBuffer1(327) <= LineBuffer1(326);
			LineBuffer1(328) <= LineBuffer1(327);
			LineBuffer1(329) <= LineBuffer1(328);	
			LineBuffer1(330) <= LineBuffer1(329);
			LineBuffer1(331) <= LineBuffer1(330);
			LineBuffer1(332) <= LineBuffer1(331);
			LineBuffer1(333) <= LineBuffer1(332);
			LineBuffer1(334) <= LineBuffer1(333);
			LineBuffer1(335) <= LineBuffer1(334);
			LineBuffer1(336) <= LineBuffer1(335);
			LineBuffer1(337) <= LineBuffer1(336);
			LineBuffer1(338) <= LineBuffer1(337);
			LineBuffer1(339) <= LineBuffer1(338);	
			LineBuffer1(340) <= LineBuffer1(339);
			LineBuffer1(341) <= LineBuffer1(340);
			LineBuffer1(342) <= LineBuffer1(341);
			LineBuffer1(343) <= LineBuffer1(342);
			LineBuffer1(344) <= LineBuffer1(343);
			LineBuffer1(345) <= LineBuffer1(344);
			LineBuffer1(346) <= LineBuffer1(345);
			LineBuffer1(347) <= LineBuffer1(346);
			LineBuffer1(348) <= LineBuffer1(347);
			LineBuffer1(349) <= LineBuffer1(348);	
			LineBuffer1(350) <= LineBuffer1(349);
			LineBuffer1(351) <= LineBuffer1(350);
			LineBuffer1(352) <= LineBuffer1(351);
			LineBuffer1(353) <= LineBuffer1(352);
			LineBuffer1(354) <= LineBuffer1(353);
			LineBuffer1(355) <= LineBuffer1(354);
			LineBuffer1(356) <= LineBuffer1(355);
			LineBuffer1(357) <= LineBuffer1(356);
			LineBuffer1(358) <= LineBuffer1(357);
			LineBuffer1(359) <= LineBuffer1(358);	
			LineBuffer1(360) <= LineBuffer1(359);
			LineBuffer1(361) <= LineBuffer1(360);
			LineBuffer1(362) <= LineBuffer1(361);
			LineBuffer1(363) <= LineBuffer1(362);
			LineBuffer1(364) <= LineBuffer1(363);
			LineBuffer1(365) <= LineBuffer1(364);
			LineBuffer1(366) <= LineBuffer1(365);
			LineBuffer1(367) <= LineBuffer1(366);
			LineBuffer1(368) <= LineBuffer1(367);
			LineBuffer1(369) <= LineBuffer1(368);	
			LineBuffer1(370) <= LineBuffer1(369);
			LineBuffer1(371) <= LineBuffer1(370);
			LineBuffer1(372) <= LineBuffer1(371);
			LineBuffer1(373) <= LineBuffer1(372);
			LineBuffer1(374) <= LineBuffer1(373);
			LineBuffer1(375) <= LineBuffer1(374);
			LineBuffer1(376) <= LineBuffer1(375);
			LineBuffer1(377) <= LineBuffer1(376);
			LineBuffer1(378) <= LineBuffer1(377);
			LineBuffer1(379) <= LineBuffer1(378);	
			LineBuffer1(380) <= LineBuffer1(379);
			LineBuffer1(381) <= LineBuffer1(380);
			LineBuffer1(382) <= LineBuffer1(381);
			LineBuffer1(383) <= LineBuffer1(382);
			LineBuffer1(384) <= LineBuffer1(383);
			LineBuffer1(385) <= LineBuffer1(384);
			LineBuffer1(386) <= LineBuffer1(385);
			LineBuffer1(387) <= LineBuffer1(386);
			LineBuffer1(388) <= LineBuffer1(387);
			LineBuffer1(389) <= LineBuffer1(388);	
			LineBuffer1(390) <= LineBuffer1(389);
			LineBuffer1(391) <= LineBuffer1(390);
			LineBuffer1(392) <= LineBuffer1(391);
			LineBuffer1(393) <= LineBuffer1(392);
			LineBuffer1(394) <= LineBuffer1(393);
			LineBuffer1(395) <= LineBuffer1(394);
			LineBuffer1(396) <= LineBuffer1(395);
			LineBuffer1(397) <= LineBuffer1(396);
			LineBuffer1(398) <= LineBuffer1(397);
			LineBuffer1(399) <= LineBuffer1(398);
			LineBuffer1(400) <= LineBuffer1(399);	
			LineBuffer1(401) <= LineBuffer1(400);
			LineBuffer1(402) <= LineBuffer1(401);
			LineBuffer1(403) <= LineBuffer1(402);
			LineBuffer1(404) <= LineBuffer1(403);
			LineBuffer1(405) <= LineBuffer1(404);
			LineBuffer1(406) <= LineBuffer1(405);
			LineBuffer1(407) <= LineBuffer1(406);
			LineBuffer1(408) <= LineBuffer1(407);
			LineBuffer1(409) <= LineBuffer1(408);	
			LineBuffer1(410) <= LineBuffer1(409);
			LineBuffer1(411) <= LineBuffer1(410);
			LineBuffer1(412) <= LineBuffer1(411);
			LineBuffer1(413) <= LineBuffer1(412);
			LineBuffer1(414) <= LineBuffer1(413);
			LineBuffer1(415) <= LineBuffer1(414);
			LineBuffer1(416) <= LineBuffer1(415);
			LineBuffer1(417) <= LineBuffer1(416);
			LineBuffer1(418) <= LineBuffer1(417);
			LineBuffer1(419) <= LineBuffer1(418);	
			LineBuffer1(420) <= LineBuffer1(419);
			LineBuffer1(421) <= LineBuffer1(420);
			LineBuffer1(422) <= LineBuffer1(421);
			LineBuffer1(423) <= LineBuffer1(422);
			LineBuffer1(424) <= LineBuffer1(423);
			LineBuffer1(425) <= LineBuffer1(424);
			LineBuffer1(426) <= LineBuffer1(425);
			LineBuffer1(427) <= LineBuffer1(426);
			LineBuffer1(428) <= LineBuffer1(427);
			LineBuffer1(429) <= LineBuffer1(428);	
			LineBuffer1(430) <= LineBuffer1(429);
			LineBuffer1(431) <= LineBuffer1(430);
			LineBuffer1(432) <= LineBuffer1(431);
			LineBuffer1(433) <= LineBuffer1(432);
			LineBuffer1(434) <= LineBuffer1(433);
			LineBuffer1(435) <= LineBuffer1(434);
			LineBuffer1(436) <= LineBuffer1(435);
			LineBuffer1(437) <= LineBuffer1(436);
			LineBuffer1(438) <= LineBuffer1(437);
			LineBuffer1(439) <= LineBuffer1(438);	
			LineBuffer1(440) <= LineBuffer1(439);
			LineBuffer1(441) <= LineBuffer1(440);
			LineBuffer1(442) <= LineBuffer1(441);
			LineBuffer1(443) <= LineBuffer1(442);
			LineBuffer1(444) <= LineBuffer1(443);
			LineBuffer1(445) <= LineBuffer1(444);
			LineBuffer1(446) <= LineBuffer1(445);
			LineBuffer1(447) <= LineBuffer1(446);
			LineBuffer1(448) <= LineBuffer1(447);
			LineBuffer1(449) <= LineBuffer1(448);	
			LineBuffer1(450) <= LineBuffer1(449);
			LineBuffer1(451) <= LineBuffer1(450);
			LineBuffer1(452) <= LineBuffer1(451);
			LineBuffer1(453) <= LineBuffer1(452);
			LineBuffer1(454) <= LineBuffer1(453);
			LineBuffer1(455) <= LineBuffer1(454);
			LineBuffer1(456) <= LineBuffer1(455);
			LineBuffer1(457) <= LineBuffer1(456);
			LineBuffer1(458) <= LineBuffer1(457);
			LineBuffer1(459) <= LineBuffer1(458);	
			LineBuffer1(460) <= LineBuffer1(459);
			LineBuffer1(461) <= LineBuffer1(460);
			LineBuffer1(462) <= LineBuffer1(461);
			LineBuffer1(463) <= LineBuffer1(462);
			LineBuffer1(464) <= LineBuffer1(463);
			LineBuffer1(465) <= LineBuffer1(464);
			LineBuffer1(466) <= LineBuffer1(465);
			LineBuffer1(467) <= LineBuffer1(466);
			LineBuffer1(468) <= LineBuffer1(467);
			LineBuffer1(469) <= LineBuffer1(468);	
			LineBuffer1(470) <= LineBuffer1(469);
			LineBuffer1(471) <= LineBuffer1(470);
			LineBuffer1(472) <= LineBuffer1(471);
			LineBuffer1(473) <= LineBuffer1(472);
			LineBuffer1(474) <= LineBuffer1(473);
			LineBuffer1(475) <= LineBuffer1(474);
			LineBuffer1(476) <= LineBuffer1(475);
			LineBuffer1(477) <= LineBuffer1(476);
			LineBuffer1(478) <= LineBuffer1(477);
			LineBuffer1(479) <= LineBuffer1(478);	
			LineBuffer1(480) <= LineBuffer1(479);
			LineBuffer1(481) <= LineBuffer1(480);
			LineBuffer1(482) <= LineBuffer1(481);
			LineBuffer1(483) <= LineBuffer1(482);
			LineBuffer1(484) <= LineBuffer1(483);
			LineBuffer1(485) <= LineBuffer1(484);
			LineBuffer1(486) <= LineBuffer1(485);
			LineBuffer1(487) <= LineBuffer1(486);
			LineBuffer1(488) <= LineBuffer1(487);
			LineBuffer1(489) <= LineBuffer1(488);	
			LineBuffer1(490) <= LineBuffer1(489);
			LineBuffer1(491) <= LineBuffer1(490);
			LineBuffer1(492) <= LineBuffer1(491);
			LineBuffer1(493) <= LineBuffer1(492);
			LineBuffer1(494) <= LineBuffer1(493);
			LineBuffer1(495) <= LineBuffer1(494);
			LineBuffer1(496) <= LineBuffer1(495);
			LineBuffer1(497) <= LineBuffer1(496);
			LineBuffer1(498) <= LineBuffer1(497);
			LineBuffer1(499) <= LineBuffer1(498);	
			LineBuffer1(500) <= LineBuffer1(499);	
			LineBuffer1(501) <= LineBuffer1(500);
			LineBuffer1(502) <= LineBuffer1(501);
			LineBuffer1(503) <= LineBuffer1(502);
			LineBuffer1(504) <= LineBuffer1(503);
			LineBuffer1(505) <= LineBuffer1(504);
			LineBuffer1(506) <= LineBuffer1(505);
			LineBuffer1(507) <= LineBuffer1(506);
			LineBuffer1(508) <= LineBuffer1(507);
			LineBuffer1(509) <= LineBuffer1(508);	
			LineBuffer1(510) <= LineBuffer1(509);
			LineBuffer1(511) <= LineBuffer1(510);
			LineBuffer1(512) <= LineBuffer1(511);
			LineBuffer1(513) <= LineBuffer1(512);
			LineBuffer1(514) <= LineBuffer1(513);
			LineBuffer1(515) <= LineBuffer1(514);
			LineBuffer1(516) <= LineBuffer1(515);
			LineBuffer1(517) <= LineBuffer1(516);
			LineBuffer1(518) <= LineBuffer1(517);
			LineBuffer1(519) <= LineBuffer1(518);	
			LineBuffer1(520) <= LineBuffer1(519);
			LineBuffer1(521) <= LineBuffer1(520);
			LineBuffer1(522) <= LineBuffer1(521);
			LineBuffer1(523) <= LineBuffer1(522);
			LineBuffer1(524) <= LineBuffer1(523);
			LineBuffer1(525) <= LineBuffer1(524);
			LineBuffer1(526) <= LineBuffer1(525);
			LineBuffer1(527) <= LineBuffer1(526);
			LineBuffer1(528) <= LineBuffer1(527);
			LineBuffer1(529) <= LineBuffer1(528);	
			LineBuffer1(530) <= LineBuffer1(529);
			LineBuffer1(531) <= LineBuffer1(530);
			LineBuffer1(532) <= LineBuffer1(531);
			LineBuffer1(533) <= LineBuffer1(532);
			LineBuffer1(534) <= LineBuffer1(533);
			LineBuffer1(535) <= LineBuffer1(534);
			LineBuffer1(536) <= LineBuffer1(535);
			LineBuffer1(537) <= LineBuffer1(536);
			LineBuffer1(538) <= LineBuffer1(537);
			LineBuffer1(539) <= LineBuffer1(538);	
			LineBuffer1(540) <= LineBuffer1(539);
			LineBuffer1(541) <= LineBuffer1(540);
			LineBuffer1(542) <= LineBuffer1(541);
			LineBuffer1(543) <= LineBuffer1(542);
			LineBuffer1(544) <= LineBuffer1(543);
			LineBuffer1(545) <= LineBuffer1(544);
			LineBuffer1(546) <= LineBuffer1(545);
			LineBuffer1(547) <= LineBuffer1(546);
			LineBuffer1(548) <= LineBuffer1(547);
			LineBuffer1(549) <= LineBuffer1(548);	
			LineBuffer1(550) <= LineBuffer1(549);
			LineBuffer1(551) <= LineBuffer1(550);
			LineBuffer1(552) <= LineBuffer1(551);
			LineBuffer1(553) <= LineBuffer1(552);
			LineBuffer1(554) <= LineBuffer1(553);
			LineBuffer1(555) <= LineBuffer1(554);
			LineBuffer1(556) <= LineBuffer1(555);
			LineBuffer1(557) <= LineBuffer1(556);
			LineBuffer1(558) <= LineBuffer1(557);
			LineBuffer1(559) <= LineBuffer1(558);	
			LineBuffer1(560) <= LineBuffer1(559);
			LineBuffer1(561) <= LineBuffer1(560);
			LineBuffer1(562) <= LineBuffer1(561);
			LineBuffer1(563) <= LineBuffer1(562);
			LineBuffer1(564) <= LineBuffer1(563);
			LineBuffer1(565) <= LineBuffer1(564);
			LineBuffer1(566) <= LineBuffer1(565);
			LineBuffer1(567) <= LineBuffer1(566);
			LineBuffer1(568) <= LineBuffer1(567);
			LineBuffer1(569) <= LineBuffer1(568);	
			LineBuffer1(570) <= LineBuffer1(569);
			LineBuffer1(571) <= LineBuffer1(570);
			LineBuffer1(572) <= LineBuffer1(571);
			LineBuffer1(573) <= LineBuffer1(572);
			LineBuffer1(574) <= LineBuffer1(573);
			LineBuffer1(575) <= LineBuffer1(574);
			LineBuffer1(576) <= LineBuffer1(575);
			LineBuffer1(577) <= LineBuffer1(576);
			LineBuffer1(578) <= LineBuffer1(577);
			LineBuffer1(579) <= LineBuffer1(578);	
			LineBuffer1(580) <= LineBuffer1(579);
			LineBuffer1(581) <= LineBuffer1(580);
			LineBuffer1(582) <= LineBuffer1(581);
			LineBuffer1(583) <= LineBuffer1(582);
			LineBuffer1(584) <= LineBuffer1(583);
			LineBuffer1(585) <= LineBuffer1(584);
			LineBuffer1(586) <= LineBuffer1(585);
			LineBuffer1(587) <= LineBuffer1(586);
			LineBuffer1(588) <= LineBuffer1(587);
			LineBuffer1(589) <= LineBuffer1(588);	
			LineBuffer1(590) <= LineBuffer1(589);
			LineBuffer1(591) <= LineBuffer1(590);
			LineBuffer1(592) <= LineBuffer1(591);
			LineBuffer1(593) <= LineBuffer1(592);
			LineBuffer1(594) <= LineBuffer1(593);
			LineBuffer1(595) <= LineBuffer1(594);
			LineBuffer1(596) <= LineBuffer1(595);
			LineBuffer1(597) <= LineBuffer1(596);
			LineBuffer1(598) <= LineBuffer1(597);
			LineBuffer1(599) <= LineBuffer1(598);	
			LineBuffer1(600) <= LineBuffer1(599);	
			LineBuffer1(601) <= LineBuffer1(600);
			LineBuffer1(602) <= LineBuffer1(601);
			LineBuffer1(603) <= LineBuffer1(602);
			LineBuffer1(604) <= LineBuffer1(603);
			LineBuffer1(605) <= LineBuffer1(604);
			LineBuffer1(606) <= LineBuffer1(605);
			LineBuffer1(607) <= LineBuffer1(606);
			LineBuffer1(608) <= LineBuffer1(607);
			LineBuffer1(609) <= LineBuffer1(608);	
			LineBuffer1(610) <= LineBuffer1(609);
			LineBuffer1(611) <= LineBuffer1(610);
			LineBuffer1(612) <= LineBuffer1(611);
			LineBuffer1(613) <= LineBuffer1(612);
			LineBuffer1(614) <= LineBuffer1(613);
			LineBuffer1(615) <= LineBuffer1(614);
			LineBuffer1(616) <= LineBuffer1(615);
			LineBuffer1(617) <= LineBuffer1(616);
			LineBuffer1(618) <= LineBuffer1(617);
			LineBuffer1(619) <= LineBuffer1(618);	
			LineBuffer1(620) <= LineBuffer1(619);
			LineBuffer1(621) <= LineBuffer1(620);
			LineBuffer1(622) <= LineBuffer1(621);
			LineBuffer1(623) <= LineBuffer1(622);
			LineBuffer1(624) <= LineBuffer1(623);
			LineBuffer1(625) <= LineBuffer1(624);
			LineBuffer1(626) <= LineBuffer1(625);
			LineBuffer1(627) <= LineBuffer1(626);
			LineBuffer1(628) <= LineBuffer1(627);
			LineBuffer1(629) <= LineBuffer1(628);	
			LineBuffer1(630) <= LineBuffer1(629);
			LineBuffer1(631) <= LineBuffer1(630);
			LineBuffer1(632) <= LineBuffer1(631);
			LineBuffer1(633) <= LineBuffer1(632);
			LineBuffer1(634) <= LineBuffer1(633);
			LineBuffer1(635) <= LineBuffer1(634);
			LineBuffer1(636) <= LineBuffer1(635);
			LineBuffer1(637) <= LineBuffer1(636);
			LineBuffer1(638) <= LineBuffer1(637);
			LineBuffer1(639) <= LineBuffer1(638);
			LineBuffer1(640) <= LineBuffer1(639);
            LineBuffer1(641) <= LineBuffer1(640);
            LineBuffer1(642) <= LineBuffer1(641);
            LineBuffer1(643) <= LineBuffer1(642);
            LineBuffer1(644) <= LineBuffer1(643);
            LineBuffer1(645) <= LineBuffer1(644);
            LineBuffer1(646) <= LineBuffer1(645);
            LineBuffer1(647) <= LineBuffer1(646);
            LineBuffer1(648) <= LineBuffer1(647);
            LineBuffer1(649) <= LineBuffer1(648);    
            LineBuffer1(650) <= LineBuffer1(649);
            LineBuffer1(651) <= LineBuffer1(650);
            LineBuffer1(652) <= LineBuffer1(651);
            LineBuffer1(653) <= LineBuffer1(652);
            LineBuffer1(654) <= LineBuffer1(653);
            LineBuffer1(655) <= LineBuffer1(654);
            LineBuffer1(656) <= LineBuffer1(655);
            LineBuffer1(657) <= LineBuffer1(656);
            LineBuffer1(658) <= LineBuffer1(657);
            LineBuffer1(659) <= LineBuffer1(658);    
            LineBuffer1(660) <= LineBuffer1(659);
            LineBuffer1(661) <= LineBuffer1(660);
            LineBuffer1(662) <= LineBuffer1(661);
            LineBuffer1(663) <= LineBuffer1(662);
            LineBuffer1(664) <= LineBuffer1(663);
            LineBuffer1(665) <= LineBuffer1(664);
            LineBuffer1(666) <= LineBuffer1(665);
            LineBuffer1(667) <= LineBuffer1(666);
            LineBuffer1(668) <= LineBuffer1(667);
            LineBuffer1(669) <= LineBuffer1(668);    
            LineBuffer1(670) <= LineBuffer1(669);
            LineBuffer1(671) <= LineBuffer1(670);
            LineBuffer1(672) <= LineBuffer1(671);
            LineBuffer1(673) <= LineBuffer1(672);
            LineBuffer1(674) <= LineBuffer1(673);
            LineBuffer1(675) <= LineBuffer1(674);
            LineBuffer1(676) <= LineBuffer1(675);
            LineBuffer1(677) <= LineBuffer1(676);
            LineBuffer1(678) <= LineBuffer1(677);
            LineBuffer1(679) <= LineBuffer1(678);    
            LineBuffer1(680) <= LineBuffer1(679);
            LineBuffer1(681) <= LineBuffer1(680);
            LineBuffer1(682) <= LineBuffer1(681);
            LineBuffer1(683) <= LineBuffer1(682);
            LineBuffer1(684) <= LineBuffer1(683);
            LineBuffer1(685) <= LineBuffer1(684);
            LineBuffer1(686) <= LineBuffer1(685);
            LineBuffer1(687) <= LineBuffer1(686);
            LineBuffer1(688) <= LineBuffer1(687);
            LineBuffer1(689) <= LineBuffer1(688);    
            LineBuffer1(690) <= LineBuffer1(689);
            LineBuffer1(691) <= LineBuffer1(690);
            LineBuffer1(692) <= LineBuffer1(691);
            LineBuffer1(693) <= LineBuffer1(692);
            LineBuffer1(694) <= LineBuffer1(693);
            LineBuffer1(695) <= LineBuffer1(694);
            LineBuffer1(696) <= LineBuffer1(695);
            LineBuffer1(697) <= LineBuffer1(696);
            LineBuffer1(698) <= LineBuffer1(697);
            LineBuffer1(699) <= LineBuffer1(698);    
            LineBuffer1(700) <= LineBuffer1(699);
            LineBuffer1(701) <= LineBuffer1(700);
            LineBuffer1(702) <= LineBuffer1(701);
            LineBuffer1(703) <= LineBuffer1(702);
            LineBuffer1(704) <= LineBuffer1(703);
            LineBuffer1(705) <= LineBuffer1(704);
            LineBuffer1(706) <= LineBuffer1(705);
            LineBuffer1(707) <= LineBuffer1(706);
            LineBuffer1(708) <= LineBuffer1(707);
            LineBuffer1(709) <= LineBuffer1(708);    
            LineBuffer1(710) <= LineBuffer1(709);
            LineBuffer1(711) <= LineBuffer1(710);
            LineBuffer1(712) <= LineBuffer1(711);
            LineBuffer1(713) <= LineBuffer1(712);
            LineBuffer1(714) <= LineBuffer1(713);
            LineBuffer1(715) <= LineBuffer1(714);
            LineBuffer1(716) <= LineBuffer1(715);
            LineBuffer1(717) <= LineBuffer1(716);
            LineBuffer1(718) <= LineBuffer1(717);
            LineBuffer1(719) <= LineBuffer1(718);    
            LineBuffer1(720) <= LineBuffer1(719);
            LineBuffer1(721) <= LineBuffer1(720);
            LineBuffer1(722) <= LineBuffer1(721);
            LineBuffer1(723) <= LineBuffer1(722);
            LineBuffer1(724) <= LineBuffer1(723);
            LineBuffer1(725) <= LineBuffer1(724);
            LineBuffer1(726) <= LineBuffer1(725);
            LineBuffer1(727) <= LineBuffer1(726);
            LineBuffer1(728) <= LineBuffer1(727);
            LineBuffer1(729) <= LineBuffer1(728);    
            LineBuffer1(730) <= LineBuffer1(729);
            LineBuffer1(731) <= LineBuffer1(730);
            LineBuffer1(732) <= LineBuffer1(731);
            LineBuffer1(733) <= LineBuffer1(732);
            LineBuffer1(734) <= LineBuffer1(733);
            LineBuffer1(735) <= LineBuffer1(734);
            LineBuffer1(736) <= LineBuffer1(735);
            LineBuffer1(737) <= LineBuffer1(736);
            LineBuffer1(738) <= LineBuffer1(737);
            LineBuffer1(739) <= LineBuffer1(738);    
            LineBuffer1(740) <= LineBuffer1(739);
            LineBuffer1(741) <= LineBuffer1(740);
            LineBuffer1(742) <= LineBuffer1(741);
            LineBuffer1(743) <= LineBuffer1(742);
            LineBuffer1(744) <= LineBuffer1(743);
            LineBuffer1(745) <= LineBuffer1(744);
            LineBuffer1(746) <= LineBuffer1(745);
            LineBuffer1(747) <= LineBuffer1(746);
            LineBuffer1(748) <= LineBuffer1(747);
            LineBuffer1(749) <= LineBuffer1(748);    
            LineBuffer1(750) <= LineBuffer1(749);
            LineBuffer1(751) <= LineBuffer1(750);
            LineBuffer1(752) <= LineBuffer1(751);
            LineBuffer1(753) <= LineBuffer1(752);
            LineBuffer1(754) <= LineBuffer1(753);
            LineBuffer1(755) <= LineBuffer1(754);
            LineBuffer1(756) <= LineBuffer1(755);
            LineBuffer1(757) <= LineBuffer1(756);
            LineBuffer1(758) <= LineBuffer1(757);
            LineBuffer1(759) <= LineBuffer1(758);    
            LineBuffer1(760) <= LineBuffer1(759);
            LineBuffer1(761) <= LineBuffer1(760);
            LineBuffer1(762) <= LineBuffer1(761);
            LineBuffer1(763) <= LineBuffer1(762);
            LineBuffer1(764) <= LineBuffer1(763);
            LineBuffer1(765) <= LineBuffer1(764);
            LineBuffer1(766) <= LineBuffer1(765);
            LineBuffer1(767) <= LineBuffer1(766);
            LineBuffer1(768) <= LineBuffer1(767);
            LineBuffer1(769) <= LineBuffer1(768);    
            LineBuffer1(770) <= LineBuffer1(769);
            LineBuffer1(771) <= LineBuffer1(770);
            LineBuffer1(772) <= LineBuffer1(771);
            LineBuffer1(773) <= LineBuffer1(772);
            LineBuffer1(774) <= LineBuffer1(773);
            LineBuffer1(775) <= LineBuffer1(774);
            LineBuffer1(776) <= LineBuffer1(775);
            LineBuffer1(777) <= LineBuffer1(776);
            LineBuffer1(778) <= LineBuffer1(777);
            LineBuffer1(779) <= LineBuffer1(778);    
            LineBuffer1(780) <= LineBuffer1(779);
            LineBuffer1(781) <= LineBuffer1(780);
            LineBuffer1(782) <= LineBuffer1(781);
            LineBuffer1(783) <= LineBuffer1(782);
            LineBuffer1(784) <= LineBuffer1(783);
            LineBuffer1(785) <= LineBuffer1(784);
            LineBuffer1(786) <= LineBuffer1(785);
            LineBuffer1(787) <= LineBuffer1(786);
            LineBuffer1(788) <= LineBuffer1(787);
            LineBuffer1(789) <= LineBuffer1(788);    
            LineBuffer1(790) <= LineBuffer1(789);
            LineBuffer1(791) <= LineBuffer1(790);
            LineBuffer1(792) <= LineBuffer1(791);
            LineBuffer1(793) <= LineBuffer1(792);
            LineBuffer1(794) <= LineBuffer1(793);
            LineBuffer1(795) <= LineBuffer1(794);
            LineBuffer1(796) <= LineBuffer1(795);
            LineBuffer1(797) <= LineBuffer1(796);
            LineBuffer1(798) <= LineBuffer1(797);
            LineBuffer1(799) <= LineBuffer1(798);    
            LineBuffer1(800) <= LineBuffer1(799);
            LineBuffer1(801) <= LineBuffer1(800);
            LineBuffer1(802) <= LineBuffer1(801);
            LineBuffer1(803) <= LineBuffer1(802);
            LineBuffer1(804) <= LineBuffer1(803);
            LineBuffer1(805) <= LineBuffer1(804);
            LineBuffer1(806) <= LineBuffer1(805);
            LineBuffer1(807) <= LineBuffer1(806);
            LineBuffer1(808) <= LineBuffer1(807);
            LineBuffer1(809) <= LineBuffer1(808);    
            LineBuffer1(810) <= LineBuffer1(809);
            LineBuffer1(811) <= LineBuffer1(810);
            LineBuffer1(812) <= LineBuffer1(811);
            LineBuffer1(813) <= LineBuffer1(812);
            LineBuffer1(814) <= LineBuffer1(813);
            LineBuffer1(815) <= LineBuffer1(814);
            LineBuffer1(816) <= LineBuffer1(815);
            LineBuffer1(817) <= LineBuffer1(816);
            LineBuffer1(818) <= LineBuffer1(817);
            LineBuffer1(819) <= LineBuffer1(818);    
            LineBuffer1(820) <= LineBuffer1(819);
            LineBuffer1(821) <= LineBuffer1(820);
            LineBuffer1(822) <= LineBuffer1(821);
            LineBuffer1(823) <= LineBuffer1(822);
            LineBuffer1(824) <= LineBuffer1(823);
            LineBuffer1(825) <= LineBuffer1(824);
            LineBuffer1(826) <= LineBuffer1(825);
            LineBuffer1(827) <= LineBuffer1(826);
            LineBuffer1(828) <= LineBuffer1(827);
            LineBuffer1(829) <= LineBuffer1(828);    
            LineBuffer1(830) <= LineBuffer1(829);
            LineBuffer1(831) <= LineBuffer1(830);
            LineBuffer1(832) <= LineBuffer1(831);
            LineBuffer1(833) <= LineBuffer1(832);
            LineBuffer1(834) <= LineBuffer1(833);
            LineBuffer1(835) <= LineBuffer1(834);
            LineBuffer1(836) <= LineBuffer1(835);
            LineBuffer1(837) <= LineBuffer1(836);
            LineBuffer1(838) <= LineBuffer1(837);
            LineBuffer1(839) <= LineBuffer1(838);
            LineBuffer1(840) <= LineBuffer1(839);
            LineBuffer1(841) <= LineBuffer1(840);
            LineBuffer1(842) <= LineBuffer1(841);
            LineBuffer1(843) <= LineBuffer1(842);
            LineBuffer1(844) <= LineBuffer1(843);
            LineBuffer1(845) <= LineBuffer1(844);
            LineBuffer1(846) <= LineBuffer1(845);
            LineBuffer1(847) <= LineBuffer1(846);
            LineBuffer1(848) <= LineBuffer1(847);
            LineBuffer1(849) <= LineBuffer1(848);    
            LineBuffer1(850) <= LineBuffer1(849);
            LineBuffer1(851) <= LineBuffer1(850);
            LineBuffer1(852) <= LineBuffer1(851);
            LineBuffer1(853) <= LineBuffer1(852);
            LineBuffer1(854) <= LineBuffer1(853);
            LineBuffer1(855) <= LineBuffer1(854);
            LineBuffer1(856) <= LineBuffer1(855);
            LineBuffer1(857) <= LineBuffer1(856);
            LineBuffer1(858) <= LineBuffer1(857);
            LineBuffer1(859) <= LineBuffer1(858);    
            LineBuffer1(860) <= LineBuffer1(859);
            LineBuffer1(861) <= LineBuffer1(860);
            LineBuffer1(862) <= LineBuffer1(861);
            LineBuffer1(863) <= LineBuffer1(862);
            LineBuffer1(864) <= LineBuffer1(863);
            LineBuffer1(865) <= LineBuffer1(864);
            LineBuffer1(866) <= LineBuffer1(865);
            LineBuffer1(867) <= LineBuffer1(866);
            LineBuffer1(868) <= LineBuffer1(867);
            LineBuffer1(869) <= LineBuffer1(868);    
            LineBuffer1(870) <= LineBuffer1(869);
            LineBuffer1(871) <= LineBuffer1(870);
            LineBuffer1(872) <= LineBuffer1(871);
            LineBuffer1(873) <= LineBuffer1(872);
            LineBuffer1(874) <= LineBuffer1(873);
            LineBuffer1(875) <= LineBuffer1(874);
            LineBuffer1(876) <= LineBuffer1(875);
            LineBuffer1(877) <= LineBuffer1(876);
            LineBuffer1(878) <= LineBuffer1(877);
            LineBuffer1(879) <= LineBuffer1(878);    
            LineBuffer1(880) <= LineBuffer1(879);
            LineBuffer1(881) <= LineBuffer1(880);
            LineBuffer1(882) <= LineBuffer1(881);
            LineBuffer1(883) <= LineBuffer1(882);
            LineBuffer1(884) <= LineBuffer1(883);
            LineBuffer1(885) <= LineBuffer1(884);
            LineBuffer1(886) <= LineBuffer1(885);
            LineBuffer1(887) <= LineBuffer1(886);
            LineBuffer1(888) <= LineBuffer1(887);
            LineBuffer1(889) <= LineBuffer1(888);    
            LineBuffer1(890) <= LineBuffer1(889);
            LineBuffer1(891) <= LineBuffer1(890);
            LineBuffer1(892) <= LineBuffer1(891);
            LineBuffer1(893) <= LineBuffer1(892);
            LineBuffer1(894) <= LineBuffer1(893);
            LineBuffer1(895) <= LineBuffer1(894);
            LineBuffer1(896) <= LineBuffer1(895);
            LineBuffer1(897) <= LineBuffer1(896);
            LineBuffer1(898) <= LineBuffer1(897);
            LineBuffer1(899) <= LineBuffer1(898);    
            LineBuffer1(900) <= LineBuffer1(899);
            LineBuffer1(901) <= LineBuffer1(900);
            LineBuffer1(902) <= LineBuffer1(901);
            LineBuffer1(903) <= LineBuffer1(902);
            LineBuffer1(904) <= LineBuffer1(903);
            LineBuffer1(905) <= LineBuffer1(904);
            LineBuffer1(906) <= LineBuffer1(905);
            LineBuffer1(907) <= LineBuffer1(906);
            LineBuffer1(908) <= LineBuffer1(907);
            LineBuffer1(909) <= LineBuffer1(908);    
            LineBuffer1(910) <= LineBuffer1(909);
            LineBuffer1(911) <= LineBuffer1(910);
            LineBuffer1(912) <= LineBuffer1(911);
            LineBuffer1(913) <= LineBuffer1(912);
            LineBuffer1(914) <= LineBuffer1(913);
            LineBuffer1(915) <= LineBuffer1(914);
            LineBuffer1(916) <= LineBuffer1(915);
            LineBuffer1(917) <= LineBuffer1(916);
            LineBuffer1(918) <= LineBuffer1(917);
            LineBuffer1(919) <= LineBuffer1(918);    
            LineBuffer1(920) <= LineBuffer1(919);
            LineBuffer1(921) <= LineBuffer1(920);
            LineBuffer1(922) <= LineBuffer1(921);
            LineBuffer1(923) <= LineBuffer1(922);
            LineBuffer1(924) <= LineBuffer1(923);
            LineBuffer1(925) <= LineBuffer1(924);
            LineBuffer1(926) <= LineBuffer1(925);
            LineBuffer1(927) <= LineBuffer1(926);
            LineBuffer1(928) <= LineBuffer1(927);
            LineBuffer1(929) <= LineBuffer1(928);    
            LineBuffer1(930) <= LineBuffer1(929);
            LineBuffer1(931) <= LineBuffer1(930);
            LineBuffer1(932) <= LineBuffer1(931);
            LineBuffer1(933) <= LineBuffer1(932);
            LineBuffer1(934) <= LineBuffer1(933);
            LineBuffer1(935) <= LineBuffer1(934);
            LineBuffer1(936) <= LineBuffer1(935);
            LineBuffer1(937) <= LineBuffer1(936);
            LineBuffer1(938) <= LineBuffer1(937);
            LineBuffer1(939) <= LineBuffer1(938);
            LineBuffer1(940) <= LineBuffer1(939);
            LineBuffer1(941) <= LineBuffer1(940);
            LineBuffer1(942) <= LineBuffer1(941);
            LineBuffer1(943) <= LineBuffer1(942);
            LineBuffer1(944) <= LineBuffer1(943);
            LineBuffer1(945) <= LineBuffer1(944);
            LineBuffer1(946) <= LineBuffer1(945);
            LineBuffer1(947) <= LineBuffer1(946);
            LineBuffer1(948) <= LineBuffer1(947);
            LineBuffer1(949) <= LineBuffer1(948);    
            LineBuffer1(950) <= LineBuffer1(949);
            LineBuffer1(951) <= LineBuffer1(950);
            LineBuffer1(952) <= LineBuffer1(951);
            LineBuffer1(953) <= LineBuffer1(952);
            LineBuffer1(954) <= LineBuffer1(953);
            LineBuffer1(955) <= LineBuffer1(954);
            LineBuffer1(956) <= LineBuffer1(955);
            LineBuffer1(957) <= LineBuffer1(956);
            LineBuffer1(958) <= LineBuffer1(957);
            LineBuffer1(959) <= LineBuffer1(958);    
            LineBuffer1(960) <= LineBuffer1(959);
            LineBuffer1(961) <= LineBuffer1(960);
            LineBuffer1(962) <= LineBuffer1(961);
            LineBuffer1(963) <= LineBuffer1(962);
            LineBuffer1(964) <= LineBuffer1(963);
            LineBuffer1(965) <= LineBuffer1(964);
            LineBuffer1(966) <= LineBuffer1(965);
            LineBuffer1(967) <= LineBuffer1(966);
            LineBuffer1(968) <= LineBuffer1(967);
            LineBuffer1(969) <= LineBuffer1(968);    
            LineBuffer1(970) <= LineBuffer1(969);
            LineBuffer1(971) <= LineBuffer1(970);
            LineBuffer1(972) <= LineBuffer1(971);
            LineBuffer1(973) <= LineBuffer1(972);
            LineBuffer1(974) <= LineBuffer1(973);
            LineBuffer1(975) <= LineBuffer1(974);
            LineBuffer1(976) <= LineBuffer1(975);
            LineBuffer1(977) <= LineBuffer1(976);
            LineBuffer1(978) <= LineBuffer1(977);
            LineBuffer1(979) <= LineBuffer1(978);    
            LineBuffer1(980) <= LineBuffer1(979);
            LineBuffer1(981) <= LineBuffer1(980);
            LineBuffer1(982) <= LineBuffer1(981);
            LineBuffer1(983) <= LineBuffer1(982);
            LineBuffer1(984) <= LineBuffer1(983);
            LineBuffer1(985) <= LineBuffer1(984);
            LineBuffer1(986) <= LineBuffer1(985);
            LineBuffer1(987) <= LineBuffer1(986);
            LineBuffer1(988) <= LineBuffer1(987);
            LineBuffer1(989) <= LineBuffer1(988);    
            LineBuffer1(990) <= LineBuffer1(989);
            LineBuffer1(991) <= LineBuffer1(990);
            LineBuffer1(992) <= LineBuffer1(991);
            LineBuffer1(993) <= LineBuffer1(992);
            LineBuffer1(994) <= LineBuffer1(993);
            LineBuffer1(995) <= LineBuffer1(994);
            LineBuffer1(996) <= LineBuffer1(995);
            LineBuffer1(997) <= LineBuffer1(996);
            LineBuffer1(998) <= LineBuffer1(997);
            LineBuffer1(999) <= LineBuffer1(998);    
            LineBuffer1(1000) <= LineBuffer1(999);
            LineBuffer1(1001) <= LineBuffer1(1000);
            LineBuffer1(1002) <= LineBuffer1(1001);
            LineBuffer1(1003) <= LineBuffer1(1002);
            LineBuffer1(1004) <= LineBuffer1(1003);
            LineBuffer1(1005) <= LineBuffer1(1004);
            LineBuffer1(1006) <= LineBuffer1(1005);
            LineBuffer1(1007) <= LineBuffer1(1006);
            LineBuffer1(1008) <= LineBuffer1(1007);
            LineBuffer1(1009) <= LineBuffer1(1008);    
            LineBuffer1(1010) <= LineBuffer1(1009);
            LineBuffer1(1011) <= LineBuffer1(1010);
            LineBuffer1(1012) <= LineBuffer1(1011);
            LineBuffer1(1013) <= LineBuffer1(1012);
            LineBuffer1(1014) <= LineBuffer1(1013);
            LineBuffer1(1015) <= LineBuffer1(1014);
            LineBuffer1(1016) <= LineBuffer1(1015);
            LineBuffer1(1017) <= LineBuffer1(1016);
            LineBuffer1(1018) <= LineBuffer1(1017);
            LineBuffer1(1019) <= LineBuffer1(1018);    
            LineBuffer1(1020) <= LineBuffer1(1019);
            LineBuffer1(1021) <= LineBuffer1(1020);
            LineBuffer1(1022) <= LineBuffer1(1021);
            LineBuffer1(1023) <= LineBuffer1(1022);
            LineBuffer1(1024) <= LineBuffer1(1023);
            LineBuffer1(1025) <= LineBuffer1(1024);
            LineBuffer1(1026) <= LineBuffer1(1025);
            LineBuffer1(1027) <= LineBuffer1(1026);
            LineBuffer1(1028) <= LineBuffer1(1027);
            LineBuffer1(1029) <= LineBuffer1(1028);    
            LineBuffer1(1030) <= LineBuffer1(1029);
            LineBuffer1(1031) <= LineBuffer1(1030);
            LineBuffer1(1032) <= LineBuffer1(1031);
            LineBuffer1(1033) <= LineBuffer1(1032);
            LineBuffer1(1034) <= LineBuffer1(1033);
            LineBuffer1(1035) <= LineBuffer1(1034);
            LineBuffer1(1036) <= LineBuffer1(1035);
            LineBuffer1(1037) <= LineBuffer1(1036);
            LineBuffer1(1038) <= LineBuffer1(1037);
            LineBuffer1(1039) <= LineBuffer1(1038);
            LineBuffer1(1040) <= LineBuffer1(1039);
            LineBuffer1(1041) <= LineBuffer1(1040);
            LineBuffer1(1042) <= LineBuffer1(1041);
            LineBuffer1(1043) <= LineBuffer1(1042);
            LineBuffer1(1044) <= LineBuffer1(1043);
            LineBuffer1(1045) <= LineBuffer1(1044);
            LineBuffer1(1046) <= LineBuffer1(1045);
            LineBuffer1(1047) <= LineBuffer1(1046);
            LineBuffer1(1048) <= LineBuffer1(1047);
            LineBuffer1(1049) <= LineBuffer1(1048);    
            LineBuffer1(1050) <= LineBuffer1(1049);
            LineBuffer1(1051) <= LineBuffer1(1050);
            LineBuffer1(1052) <= LineBuffer1(1051);
            LineBuffer1(1053) <= LineBuffer1(1052);
            LineBuffer1(1054) <= LineBuffer1(1053);
            LineBuffer1(1055) <= LineBuffer1(1054);
            LineBuffer1(1056) <= LineBuffer1(1055);
            LineBuffer1(1057) <= LineBuffer1(1056);
            LineBuffer1(1058) <= LineBuffer1(1057);
            LineBuffer1(1059) <= LineBuffer1(1058);    
            LineBuffer1(1060) <= LineBuffer1(1059);
            LineBuffer1(1061) <= LineBuffer1(1060);
            LineBuffer1(1062) <= LineBuffer1(1061);
            LineBuffer1(1063) <= LineBuffer1(1062);
            LineBuffer1(1064) <= LineBuffer1(1063);
            LineBuffer1(1065) <= LineBuffer1(1064);
            LineBuffer1(1066) <= LineBuffer1(1065);
            LineBuffer1(1067) <= LineBuffer1(1066);
            LineBuffer1(1068) <= LineBuffer1(1067);
            LineBuffer1(1069) <= LineBuffer1(1068);    
            LineBuffer1(1070) <= LineBuffer1(1069);
            LineBuffer1(1071) <= LineBuffer1(1070);
            LineBuffer1(1072) <= LineBuffer1(1071);
            LineBuffer1(1073) <= LineBuffer1(1072);
            LineBuffer1(1074) <= LineBuffer1(1073);
            LineBuffer1(1075) <= LineBuffer1(1074);
            LineBuffer1(1076) <= LineBuffer1(1075);
            LineBuffer1(1077) <= LineBuffer1(1076);
            LineBuffer1(1078) <= LineBuffer1(1077);
            LineBuffer1(1079) <= LineBuffer1(1078);    
            LineBuffer1(1080) <= LineBuffer1(1079);
            LineBuffer1(1081) <= LineBuffer1(1080);
            LineBuffer1(1082) <= LineBuffer1(1081);
            LineBuffer1(1083) <= LineBuffer1(1082);
            LineBuffer1(1084) <= LineBuffer1(1083);
            LineBuffer1(1085) <= LineBuffer1(1084);
            LineBuffer1(1086) <= LineBuffer1(1085);
            LineBuffer1(1087) <= LineBuffer1(1086);
            LineBuffer1(1088) <= LineBuffer1(1087);
            LineBuffer1(1089) <= LineBuffer1(1088);    
            LineBuffer1(1090) <= LineBuffer1(1089);
            LineBuffer1(1091) <= LineBuffer1(1090);
            LineBuffer1(1092) <= LineBuffer1(1091);
            LineBuffer1(1093) <= LineBuffer1(1092);
            LineBuffer1(1094) <= LineBuffer1(1093);
            LineBuffer1(1095) <= LineBuffer1(1094);
            LineBuffer1(1096) <= LineBuffer1(1095);
            LineBuffer1(1097) <= LineBuffer1(1096);
            LineBuffer1(1098) <= LineBuffer1(1097);
            LineBuffer1(1099) <= LineBuffer1(1098);    
            LineBuffer1(1100) <= LineBuffer1(1099);
            LineBuffer1(1101) <= LineBuffer1(1100);
            LineBuffer1(1102) <= LineBuffer1(1101);
            LineBuffer1(1103) <= LineBuffer1(1102);
            LineBuffer1(1104) <= LineBuffer1(1103);
            LineBuffer1(1105) <= LineBuffer1(1104);
            LineBuffer1(1106) <= LineBuffer1(1105);
            LineBuffer1(1107) <= LineBuffer1(1106);
            LineBuffer1(1108) <= LineBuffer1(1107);
            LineBuffer1(1109) <= LineBuffer1(1108);    
            LineBuffer1(1110) <= LineBuffer1(1109);
            LineBuffer1(1111) <= LineBuffer1(1110);
            LineBuffer1(1112) <= LineBuffer1(1111);
            LineBuffer1(1113) <= LineBuffer1(1112);
            LineBuffer1(1114) <= LineBuffer1(1113);
            LineBuffer1(1115) <= LineBuffer1(1114);
            LineBuffer1(1116) <= LineBuffer1(1115);
            LineBuffer1(1117) <= LineBuffer1(1116);
            LineBuffer1(1118) <= LineBuffer1(1117);
            LineBuffer1(1119) <= LineBuffer1(1118);    
            LineBuffer1(1120) <= LineBuffer1(1119);
            LineBuffer1(1121) <= LineBuffer1(1120);
            LineBuffer1(1122) <= LineBuffer1(1121);
            LineBuffer1(1123) <= LineBuffer1(1122);
            LineBuffer1(1124) <= LineBuffer1(1123);
            LineBuffer1(1125) <= LineBuffer1(1124);
            LineBuffer1(1126) <= LineBuffer1(1125);
            LineBuffer1(1127) <= LineBuffer1(1126);
            LineBuffer1(1128) <= LineBuffer1(1127);
            LineBuffer1(1129) <= LineBuffer1(1128);    
            LineBuffer1(1130) <= LineBuffer1(1129);
            LineBuffer1(1131) <= LineBuffer1(1130);
            LineBuffer1(1132) <= LineBuffer1(1131);
            LineBuffer1(1133) <= LineBuffer1(1132);
            LineBuffer1(1134) <= LineBuffer1(1133);
            LineBuffer1(1135) <= LineBuffer1(1134);
            LineBuffer1(1136) <= LineBuffer1(1135);
            LineBuffer1(1137) <= LineBuffer1(1136);
            LineBuffer1(1138) <= LineBuffer1(1137);
            LineBuffer1(1139) <= LineBuffer1(1138);
            LineBuffer1(1140) <= LineBuffer1(1139);
            LineBuffer1(1141) <= LineBuffer1(1140);
            LineBuffer1(1142) <= LineBuffer1(1141);
            LineBuffer1(1143) <= LineBuffer1(1142);
            LineBuffer1(1144) <= LineBuffer1(1143);
            LineBuffer1(1145) <= LineBuffer1(1144);
            LineBuffer1(1146) <= LineBuffer1(1145);
            LineBuffer1(1147) <= LineBuffer1(1146);
            LineBuffer1(1148) <= LineBuffer1(1147);
            LineBuffer1(1149) <= LineBuffer1(1148);    
            LineBuffer1(1150) <= LineBuffer1(1149);
            LineBuffer1(1151) <= LineBuffer1(1150);
            LineBuffer1(1152) <= LineBuffer1(1151);
            LineBuffer1(1153) <= LineBuffer1(1152);
            LineBuffer1(1154) <= LineBuffer1(1153);
            LineBuffer1(1155) <= LineBuffer1(1154);
            LineBuffer1(1156) <= LineBuffer1(1155);
            LineBuffer1(1157) <= LineBuffer1(1156);
            LineBuffer1(1158) <= LineBuffer1(1157);
            LineBuffer1(1159) <= LineBuffer1(1158);    
            LineBuffer1(1160) <= LineBuffer1(1159);
            LineBuffer1(1161) <= LineBuffer1(1160);
            LineBuffer1(1162) <= LineBuffer1(1161);
            LineBuffer1(1163) <= LineBuffer1(1162);
            LineBuffer1(1164) <= LineBuffer1(1163);
            LineBuffer1(1165) <= LineBuffer1(1164);
            LineBuffer1(1166) <= LineBuffer1(1165);
            LineBuffer1(1167) <= LineBuffer1(1166);
            LineBuffer1(1168) <= LineBuffer1(1167);
            LineBuffer1(1169) <= LineBuffer1(1168);    
            LineBuffer1(1170) <= LineBuffer1(1169);
            LineBuffer1(1171) <= LineBuffer1(1170);
            LineBuffer1(1172) <= LineBuffer1(1171);
            LineBuffer1(1173) <= LineBuffer1(1172);
            LineBuffer1(1174) <= LineBuffer1(1173);
            LineBuffer1(1175) <= LineBuffer1(1174);
            LineBuffer1(1176) <= LineBuffer1(1175);
            LineBuffer1(1177) <= LineBuffer1(1176);
            LineBuffer1(1178) <= LineBuffer1(1177);
            LineBuffer1(1179) <= LineBuffer1(1178);    
            LineBuffer1(1180) <= LineBuffer1(1179);
            LineBuffer1(1181) <= LineBuffer1(1180);
            LineBuffer1(1182) <= LineBuffer1(1181);
            LineBuffer1(1183) <= LineBuffer1(1182);
            LineBuffer1(1184) <= LineBuffer1(1183);
            LineBuffer1(1185) <= LineBuffer1(1184);
            LineBuffer1(1186) <= LineBuffer1(1185);
            LineBuffer1(1187) <= LineBuffer1(1186);
            LineBuffer1(1188) <= LineBuffer1(1187);
            LineBuffer1(1189) <= LineBuffer1(1188);    
            LineBuffer1(1190) <= LineBuffer1(1189);
            LineBuffer1(1191) <= LineBuffer1(1190);
            LineBuffer1(1192) <= LineBuffer1(1191);
            LineBuffer1(1193) <= LineBuffer1(1192);
            LineBuffer1(1194) <= LineBuffer1(1193);
            LineBuffer1(1195) <= LineBuffer1(1194);
            LineBuffer1(1196) <= LineBuffer1(1195);
            LineBuffer1(1197) <= LineBuffer1(1196);
            LineBuffer1(1198) <= LineBuffer1(1197);
            LineBuffer1(1199) <= LineBuffer1(1198);    
            LineBuffer1(1200) <= LineBuffer1(1199);
            LineBuffer1(1201) <= LineBuffer1(1200);
            LineBuffer1(1202) <= LineBuffer1(1201);
            LineBuffer1(1203) <= LineBuffer1(1202);
            LineBuffer1(1204) <= LineBuffer1(1203);
            LineBuffer1(1205) <= LineBuffer1(1204);
            LineBuffer1(1206) <= LineBuffer1(1205);
            LineBuffer1(1207) <= LineBuffer1(1206);
            LineBuffer1(1208) <= LineBuffer1(1207);
            LineBuffer1(1209) <= LineBuffer1(1208);    
            LineBuffer1(1210) <= LineBuffer1(1209);
            LineBuffer1(1211) <= LineBuffer1(1210);
            LineBuffer1(1212) <= LineBuffer1(1211);
            LineBuffer1(1213) <= LineBuffer1(1212);
            LineBuffer1(1214) <= LineBuffer1(1213);
            LineBuffer1(1215) <= LineBuffer1(1214);
            LineBuffer1(1216) <= LineBuffer1(1215);
            LineBuffer1(1217) <= LineBuffer1(1216);
            LineBuffer1(1218) <= LineBuffer1(1217);
            LineBuffer1(1219) <= LineBuffer1(1218);    
            LineBuffer1(1220) <= LineBuffer1(1219);
            LineBuffer1(1221) <= LineBuffer1(1220);
            LineBuffer1(1222) <= LineBuffer1(1221);
            LineBuffer1(1223) <= LineBuffer1(1222);
            LineBuffer1(1224) <= LineBuffer1(1223);
            LineBuffer1(1225) <= LineBuffer1(1224);
            LineBuffer1(1226) <= LineBuffer1(1225);
            LineBuffer1(1227) <= LineBuffer1(1226);
            LineBuffer1(1228) <= LineBuffer1(1227);
            LineBuffer1(1229) <= LineBuffer1(1228);    
            LineBuffer1(1230) <= LineBuffer1(1229);
            LineBuffer1(1231) <= LineBuffer1(1230);
            LineBuffer1(1232) <= LineBuffer1(1231);
            LineBuffer1(1233) <= LineBuffer1(1232);
            LineBuffer1(1234) <= LineBuffer1(1233);
            LineBuffer1(1235) <= LineBuffer1(1234);
            LineBuffer1(1236) <= LineBuffer1(1235);
            LineBuffer1(1237) <= LineBuffer1(1236);
            LineBuffer1(1238) <= LineBuffer1(1237);
            LineBuffer1(1239) <= LineBuffer1(1238);
            LineBuffer1(1240) <= LineBuffer1(1239);
            LineBuffer1(1241) <= LineBuffer1(1240);
            LineBuffer1(1242) <= LineBuffer1(1241);
            LineBuffer1(1243) <= LineBuffer1(1242);
            LineBuffer1(1244) <= LineBuffer1(1243);
            LineBuffer1(1245) <= LineBuffer1(1244);
            LineBuffer1(1246) <= LineBuffer1(1245);
            LineBuffer1(1247) <= LineBuffer1(1246);
            LineBuffer1(1248) <= LineBuffer1(1247);
            LineBuffer1(1249) <= LineBuffer1(1248);    
            LineBuffer1(1250) <= LineBuffer1(1249);
            LineBuffer1(1251) <= LineBuffer1(1250);
            LineBuffer1(1252) <= LineBuffer1(1251);
            LineBuffer1(1253) <= LineBuffer1(1252);
            LineBuffer1(1254) <= LineBuffer1(1253);
            LineBuffer1(1255) <= LineBuffer1(1254);
            LineBuffer1(1256) <= LineBuffer1(1255);
            LineBuffer1(1257) <= LineBuffer1(1256);
            LineBuffer1(1258) <= LineBuffer1(1257);
            LineBuffer1(1259) <= LineBuffer1(1258);    
            LineBuffer1(1260) <= LineBuffer1(1259);
            LineBuffer1(1261) <= LineBuffer1(1260);
            LineBuffer1(1262) <= LineBuffer1(1261);
            LineBuffer1(1263) <= LineBuffer1(1262);
            LineBuffer1(1264) <= LineBuffer1(1263);
            LineBuffer1(1265) <= LineBuffer1(1264);
            LineBuffer1(1266) <= LineBuffer1(1265);
            LineBuffer1(1267) <= LineBuffer1(1266);
            LineBuffer1(1268) <= LineBuffer1(1267);
            LineBuffer1(1269) <= LineBuffer1(1268);    
            LineBuffer1(1270) <= LineBuffer1(1269);
            LineBuffer1(1271) <= LineBuffer1(1270);
            LineBuffer1(1272) <= LineBuffer1(1271);
            LineBuffer1(1273) <= LineBuffer1(1272);
            LineBuffer1(1274) <= LineBuffer1(1273);
            LineBuffer1(1275) <= LineBuffer1(1274);
            LineBuffer1(1276) <= LineBuffer1(1275);
            LineBuffer1(1277) <= LineBuffer1(1276);
            LineBuffer1(1278) <= LineBuffer1(1277);
            LineBuffer1(1279) <= LineBuffer1(1278);
--            LineBuffer1(1280) <= LineBuffer1(1279);
--            LineBuffer1(1281) <= LineBuffer1(1280);
--            LineBuffer1(1282) <= LineBuffer1(1281);
--            LineBuffer1(1283) <= LineBuffer1(1282);
--            LineBuffer1(1284) <= LineBuffer1(1283);
--            LineBuffer1(1285) <= LineBuffer1(1284);
--            LineBuffer1(1286) <= LineBuffer1(1285);
--            LineBuffer1(1287) <= LineBuffer1(1286);
--            LineBuffer1(1288) <= LineBuffer1(1287);
--            LineBuffer1(1289) <= LineBuffer1(1288);    
--            LineBuffer1(1290) <= LineBuffer1(1289);
--            LineBuffer1(1291) <= LineBuffer1(1290);
--            LineBuffer1(1292) <= LineBuffer1(1291);
--            LineBuffer1(1293) <= LineBuffer1(1292);
--            LineBuffer1(1294) <= LineBuffer1(1293);
--            LineBuffer1(1295) <= LineBuffer1(1294);
--            LineBuffer1(1296) <= LineBuffer1(1295);
--            LineBuffer1(1297) <= LineBuffer1(1296);
--            LineBuffer1(1298) <= LineBuffer1(1297);
--            LineBuffer1(1299) <= LineBuffer1(1298);    
--            LineBuffer1(1300) <= LineBuffer1(1299);
--            LineBuffer1(1301) <= LineBuffer1(1300);
--            LineBuffer1(1302) <= LineBuffer1(1301);
--            LineBuffer1(1303) <= LineBuffer1(1302);
--            LineBuffer1(1304) <= LineBuffer1(1303);
--            LineBuffer1(1305) <= LineBuffer1(1304);
--            LineBuffer1(1306) <= LineBuffer1(1305);
--            LineBuffer1(1307) <= LineBuffer1(1306);
--            LineBuffer1(1308) <= LineBuffer1(1307);
--            LineBuffer1(1309) <= LineBuffer1(1308);    
--            LineBuffer1(1310) <= LineBuffer1(1309);
--            LineBuffer1(1311) <= LineBuffer1(1310);
--            LineBuffer1(1312) <= LineBuffer1(1311);
--            LineBuffer1(1313) <= LineBuffer1(1312);
--            LineBuffer1(1314) <= LineBuffer1(1313);
--            LineBuffer1(1315) <= LineBuffer1(1314);
--            LineBuffer1(1316) <= LineBuffer1(1315);
--            LineBuffer1(1317) <= LineBuffer1(1316);
--            LineBuffer1(1318) <= LineBuffer1(1317);
--            LineBuffer1(1319) <= LineBuffer1(1318);    
--            LineBuffer1(1320) <= LineBuffer1(1319);
--            LineBuffer1(1321) <= LineBuffer1(1320);
--            LineBuffer1(1322) <= LineBuffer1(1321);
--            LineBuffer1(1323) <= LineBuffer1(1322);
--            LineBuffer1(1324) <= LineBuffer1(1323);
--            LineBuffer1(1325) <= LineBuffer1(1324);
--            LineBuffer1(1326) <= LineBuffer1(1325);
--            LineBuffer1(1327) <= LineBuffer1(1326);
--            LineBuffer1(1328) <= LineBuffer1(1327);
--            LineBuffer1(1329) <= LineBuffer1(1328);    
--            LineBuffer1(1330) <= LineBuffer1(1329);
--            LineBuffer1(1331) <= LineBuffer1(1330);
--            LineBuffer1(1332) <= LineBuffer1(1331);
--            LineBuffer1(1333) <= LineBuffer1(1332);
--            LineBuffer1(1334) <= LineBuffer1(1333);
--            LineBuffer1(1335) <= LineBuffer1(1334);
--            LineBuffer1(1336) <= LineBuffer1(1335);
--            LineBuffer1(1337) <= LineBuffer1(1336);
--            LineBuffer1(1338) <= LineBuffer1(1337);
--            LineBuffer1(1339) <= LineBuffer1(1338);    
--            LineBuffer1(1340) <= LineBuffer1(1339);
--            LineBuffer1(1341) <= LineBuffer1(1340);
--            LineBuffer1(1342) <= LineBuffer1(1341);
--            LineBuffer1(1343) <= LineBuffer1(1342);
--            LineBuffer1(1344) <= LineBuffer1(1343);
--            LineBuffer1(1345) <= LineBuffer1(1344);
--            LineBuffer1(1346) <= LineBuffer1(1345);
--            LineBuffer1(1347) <= LineBuffer1(1346);
--            LineBuffer1(1348) <= LineBuffer1(1347);
--            LineBuffer1(1349) <= LineBuffer1(1348);    
--            LineBuffer1(1350) <= LineBuffer1(1349);
--            LineBuffer1(1351) <= LineBuffer1(1350);
--            LineBuffer1(1352) <= LineBuffer1(1351);
--            LineBuffer1(1353) <= LineBuffer1(1352);
--            LineBuffer1(1354) <= LineBuffer1(1353);
--            LineBuffer1(1355) <= LineBuffer1(1354);
--            LineBuffer1(1356) <= LineBuffer1(1355);
--            LineBuffer1(1357) <= LineBuffer1(1356);
--            LineBuffer1(1358) <= LineBuffer1(1357);
--            LineBuffer1(1359) <= LineBuffer1(1358);    
--            LineBuffer1(1360) <= LineBuffer1(1359);
--            LineBuffer1(1361) <= LineBuffer1(1360);
--            LineBuffer1(1362) <= LineBuffer1(1361);
--            LineBuffer1(1363) <= LineBuffer1(1362);
--            LineBuffer1(1364) <= LineBuffer1(1363);
--            LineBuffer1(1365) <= LineBuffer1(1364);
--            LineBuffer1(1366) <= LineBuffer1(1365);
--            LineBuffer1(1367) <= LineBuffer1(1366);
--            LineBuffer1(1368) <= LineBuffer1(1367);
--            LineBuffer1(1369) <= LineBuffer1(1368);    
--            LineBuffer1(1370) <= LineBuffer1(1369);
--            LineBuffer1(1371) <= LineBuffer1(1370);
--            LineBuffer1(1372) <= LineBuffer1(1371);
--            LineBuffer1(1373) <= LineBuffer1(1372);
--            LineBuffer1(1374) <= LineBuffer1(1373);
--            LineBuffer1(1375) <= LineBuffer1(1374);
--            LineBuffer1(1376) <= LineBuffer1(1375);
--            LineBuffer1(1377) <= LineBuffer1(1376);
--            LineBuffer1(1378) <= LineBuffer1(1377);
--            LineBuffer1(1379) <= LineBuffer1(1378);    
--            LineBuffer1(1380) <= LineBuffer1(1379);
--            LineBuffer1(1381) <= LineBuffer1(1380);
--            LineBuffer1(1382) <= LineBuffer1(1381);
--            LineBuffer1(1383) <= LineBuffer1(1382);
--            LineBuffer1(1384) <= LineBuffer1(1383);
--            LineBuffer1(1385) <= LineBuffer1(1384);
--            LineBuffer1(1386) <= LineBuffer1(1385);
--            LineBuffer1(1387) <= LineBuffer1(1386);
--            LineBuffer1(1388) <= LineBuffer1(1387);
--            LineBuffer1(1389) <= LineBuffer1(1388);    
--            LineBuffer1(1390) <= LineBuffer1(1389);
--            LineBuffer1(1391) <= LineBuffer1(1390);
--            LineBuffer1(1392) <= LineBuffer1(1391);
--            LineBuffer1(1393) <= LineBuffer1(1392);
--            LineBuffer1(1394) <= LineBuffer1(1393);
--            LineBuffer1(1395) <= LineBuffer1(1394);
--            LineBuffer1(1396) <= LineBuffer1(1395);
--            LineBuffer1(1397) <= LineBuffer1(1396);
--            LineBuffer1(1398) <= LineBuffer1(1397);
--            LineBuffer1(1399) <= LineBuffer1(1398);    
--            LineBuffer1(1400) <= LineBuffer1(1399);
--            LineBuffer1(1401) <= LineBuffer1(1400);
--            LineBuffer1(1402) <= LineBuffer1(1401);
--            LineBuffer1(1403) <= LineBuffer1(1402);
--            LineBuffer1(1404) <= LineBuffer1(1403);
--            LineBuffer1(1405) <= LineBuffer1(1404);
--            LineBuffer1(1406) <= LineBuffer1(1405);
--            LineBuffer1(1407) <= LineBuffer1(1406);
--            LineBuffer1(1408) <= LineBuffer1(1407);
--            LineBuffer1(1409) <= LineBuffer1(1408);    
--            LineBuffer1(1410) <= LineBuffer1(1409);
--            LineBuffer1(1411) <= LineBuffer1(1410);
--            LineBuffer1(1412) <= LineBuffer1(1411);
--            LineBuffer1(1413) <= LineBuffer1(1412);
--            LineBuffer1(1414) <= LineBuffer1(1413);
--            LineBuffer1(1415) <= LineBuffer1(1414);
--            LineBuffer1(1416) <= LineBuffer1(1415);
--            LineBuffer1(1417) <= LineBuffer1(1416);
--            LineBuffer1(1418) <= LineBuffer1(1417);
--            LineBuffer1(1419) <= LineBuffer1(1418);    
--            LineBuffer1(1420) <= LineBuffer1(1419);
--            LineBuffer1(1421) <= LineBuffer1(1420);
--            LineBuffer1(1422) <= LineBuffer1(1421);
--            LineBuffer1(1423) <= LineBuffer1(1422);
--            LineBuffer1(1424) <= LineBuffer1(1423);
--            LineBuffer1(1425) <= LineBuffer1(1424);
--            LineBuffer1(1426) <= LineBuffer1(1425);
--            LineBuffer1(1427) <= LineBuffer1(1426);
--            LineBuffer1(1428) <= LineBuffer1(1427);
--            LineBuffer1(1429) <= LineBuffer1(1428);    
--            LineBuffer1(1430) <= LineBuffer1(1429);
--            LineBuffer1(1431) <= LineBuffer1(1430);
--            LineBuffer1(1432) <= LineBuffer1(1431);
--            LineBuffer1(1433) <= LineBuffer1(1432);
--            LineBuffer1(1434) <= LineBuffer1(1433);
--            LineBuffer1(1435) <= LineBuffer1(1434);
--            LineBuffer1(1436) <= LineBuffer1(1435);
--            LineBuffer1(1437) <= LineBuffer1(1436);
--            LineBuffer1(1438) <= LineBuffer1(1437);
--            LineBuffer1(1439) <= LineBuffer1(1438);    
--            LineBuffer1(1440) <= LineBuffer1(1439);
--            LineBuffer1(1441) <= LineBuffer1(1440);
--            LineBuffer1(1442) <= LineBuffer1(1441);
--            LineBuffer1(1443) <= LineBuffer1(1442);
--            LineBuffer1(1444) <= LineBuffer1(1443);
--            LineBuffer1(1445) <= LineBuffer1(1444);
--            LineBuffer1(1446) <= LineBuffer1(1445);
--            LineBuffer1(1447) <= LineBuffer1(1446);
--            LineBuffer1(1448) <= LineBuffer1(1447);
--            LineBuffer1(1449) <= LineBuffer1(1448);    
--            LineBuffer1(1450) <= LineBuffer1(1449);
--            LineBuffer1(1451) <= LineBuffer1(1450);
--            LineBuffer1(1452) <= LineBuffer1(1451);
--            LineBuffer1(1453) <= LineBuffer1(1452);
--            LineBuffer1(1454) <= LineBuffer1(1453);
--            LineBuffer1(1455) <= LineBuffer1(1454);
--            LineBuffer1(1456) <= LineBuffer1(1455);
--            LineBuffer1(1457) <= LineBuffer1(1456);
--            LineBuffer1(1458) <= LineBuffer1(1457);
--            LineBuffer1(1459) <= LineBuffer1(1458);    
--            LineBuffer1(1460) <= LineBuffer1(1459);
--            LineBuffer1(1461) <= LineBuffer1(1460);
--            LineBuffer1(1462) <= LineBuffer1(1461);
--            LineBuffer1(1463) <= LineBuffer1(1462);
--            LineBuffer1(1464) <= LineBuffer1(1463);
--            LineBuffer1(1465) <= LineBuffer1(1464);
--            LineBuffer1(1466) <= LineBuffer1(1465);
--            LineBuffer1(1467) <= LineBuffer1(1466);
--            LineBuffer1(1468) <= LineBuffer1(1467);
--            LineBuffer1(1469) <= LineBuffer1(1468);    
--            LineBuffer1(1470) <= LineBuffer1(1469);
--            LineBuffer1(1471) <= LineBuffer1(1470);
--            LineBuffer1(1472) <= LineBuffer1(1471);
--            LineBuffer1(1473) <= LineBuffer1(1472);
--            LineBuffer1(1474) <= LineBuffer1(1473);
--            LineBuffer1(1475) <= LineBuffer1(1474);
--            LineBuffer1(1476) <= LineBuffer1(1475);
--            LineBuffer1(1477) <= LineBuffer1(1476);
--            LineBuffer1(1478) <= LineBuffer1(1477);
--            LineBuffer1(1479) <= LineBuffer1(1478);
--            LineBuffer1(1480) <= LineBuffer1(1479);
--            LineBuffer1(1481) <= LineBuffer1(1480);
--            LineBuffer1(1482) <= LineBuffer1(1481);
--            LineBuffer1(1483) <= LineBuffer1(1482);
--            LineBuffer1(1484) <= LineBuffer1(1483);
--            LineBuffer1(1485) <= LineBuffer1(1484);
--            LineBuffer1(1486) <= LineBuffer1(1485);
--            LineBuffer1(1487) <= LineBuffer1(1486);
--            LineBuffer1(1488) <= LineBuffer1(1487);
--            LineBuffer1(1489) <= LineBuffer1(1488);    
--            LineBuffer1(1490) <= LineBuffer1(1489);
--            LineBuffer1(1491) <= LineBuffer1(1490);
--            LineBuffer1(1492) <= LineBuffer1(1491);
--            LineBuffer1(1493) <= LineBuffer1(1492);
--            LineBuffer1(1494) <= LineBuffer1(1493);
--            LineBuffer1(1495) <= LineBuffer1(1494);
--            LineBuffer1(1496) <= LineBuffer1(1495);
--            LineBuffer1(1497) <= LineBuffer1(1496);
--            LineBuffer1(1498) <= LineBuffer1(1497);
--            LineBuffer1(1499) <= LineBuffer1(1498);    
--            LineBuffer1(1500) <= LineBuffer1(1499);
--            LineBuffer1(1501) <= LineBuffer1(1500);
--            LineBuffer1(1502) <= LineBuffer1(1501);
--            LineBuffer1(1503) <= LineBuffer1(1502);
--            LineBuffer1(1504) <= LineBuffer1(1503);
--            LineBuffer1(1505) <= LineBuffer1(1504);
--            LineBuffer1(1506) <= LineBuffer1(1505);
--            LineBuffer1(1507) <= LineBuffer1(1506);
--            LineBuffer1(1508) <= LineBuffer1(1507);
--            LineBuffer1(1509) <= LineBuffer1(1508);    
--            LineBuffer1(1510) <= LineBuffer1(1509);
--            LineBuffer1(1511) <= LineBuffer1(1510);
--            LineBuffer1(1512) <= LineBuffer1(1511);
--            LineBuffer1(1513) <= LineBuffer1(1512);
--            LineBuffer1(1514) <= LineBuffer1(1513);
--            LineBuffer1(1515) <= LineBuffer1(1514);
--            LineBuffer1(1516) <= LineBuffer1(1515);
--            LineBuffer1(1517) <= LineBuffer1(1516);
--            LineBuffer1(1518) <= LineBuffer1(1517);
--            LineBuffer1(1519) <= LineBuffer1(1518);    
--            LineBuffer1(1520) <= LineBuffer1(1519);
--            LineBuffer1(1521) <= LineBuffer1(1520);
--            LineBuffer1(1522) <= LineBuffer1(1521);
--            LineBuffer1(1523) <= LineBuffer1(1522);
--            LineBuffer1(1524) <= LineBuffer1(1523);
--            LineBuffer1(1525) <= LineBuffer1(1524);
--            LineBuffer1(1526) <= LineBuffer1(1525);
--            LineBuffer1(1527) <= LineBuffer1(1526);
--            LineBuffer1(1528) <= LineBuffer1(1527);
--            LineBuffer1(1529) <= LineBuffer1(1528);    
--            LineBuffer1(1530) <= LineBuffer1(1529);
--            LineBuffer1(1531) <= LineBuffer1(1530);
--            LineBuffer1(1532) <= LineBuffer1(1531);
--            LineBuffer1(1533) <= LineBuffer1(1532);
--            LineBuffer1(1534) <= LineBuffer1(1533);
--            LineBuffer1(1535) <= LineBuffer1(1534);
--            LineBuffer1(1536) <= LineBuffer1(1535);
--            LineBuffer1(1537) <= LineBuffer1(1536);
--            LineBuffer1(1538) <= LineBuffer1(1537);
--            LineBuffer1(1539) <= LineBuffer1(1538);    
--            LineBuffer1(1540) <= LineBuffer1(1539);
--            LineBuffer1(1541) <= LineBuffer1(1540);
--            LineBuffer1(1542) <= LineBuffer1(1541);
--            LineBuffer1(1543) <= LineBuffer1(1542);
--            LineBuffer1(1544) <= LineBuffer1(1543);
--            LineBuffer1(1545) <= LineBuffer1(1544);
--            LineBuffer1(1546) <= LineBuffer1(1545);
--            LineBuffer1(1547) <= LineBuffer1(1546);
--            LineBuffer1(1548) <= LineBuffer1(1547);
--            LineBuffer1(1549) <= LineBuffer1(1548);    
--            LineBuffer1(1550) <= LineBuffer1(1549);
--            LineBuffer1(1551) <= LineBuffer1(1550);
--            LineBuffer1(1552) <= LineBuffer1(1551);
--            LineBuffer1(1553) <= LineBuffer1(1552);
--            LineBuffer1(1554) <= LineBuffer1(1553);
--            LineBuffer1(1555) <= LineBuffer1(1554);
--            LineBuffer1(1556) <= LineBuffer1(1555);
--            LineBuffer1(1557) <= LineBuffer1(1556);
--            LineBuffer1(1558) <= LineBuffer1(1557);
--            LineBuffer1(1559) <= LineBuffer1(1558);    
--            LineBuffer1(1560) <= LineBuffer1(1559);
--            LineBuffer1(1561) <= LineBuffer1(1560);
--            LineBuffer1(1562) <= LineBuffer1(1561);
--            LineBuffer1(1563) <= LineBuffer1(1562);
--            LineBuffer1(1564) <= LineBuffer1(1563);
--            LineBuffer1(1565) <= LineBuffer1(1564);
--            LineBuffer1(1566) <= LineBuffer1(1565);
--            LineBuffer1(1567) <= LineBuffer1(1566);
--            LineBuffer1(1568) <= LineBuffer1(1567);
--            LineBuffer1(1569) <= LineBuffer1(1568);    
--            LineBuffer1(1570) <= LineBuffer1(1569);
--            LineBuffer1(1571) <= LineBuffer1(1570);
--            LineBuffer1(1572) <= LineBuffer1(1571);
--            LineBuffer1(1573) <= LineBuffer1(1572);
--            LineBuffer1(1574) <= LineBuffer1(1573);
--            LineBuffer1(1575) <= LineBuffer1(1574);
--            LineBuffer1(1576) <= LineBuffer1(1575);
--            LineBuffer1(1577) <= LineBuffer1(1576);
--            LineBuffer1(1578) <= LineBuffer1(1577);
--            LineBuffer1(1579) <= LineBuffer1(1578);
--            LineBuffer1(1580) <= LineBuffer1(1579);
--            LineBuffer1(1581) <= LineBuffer1(1580);
--            LineBuffer1(1582) <= LineBuffer1(1581);
--            LineBuffer1(1583) <= LineBuffer1(1582);
--            LineBuffer1(1584) <= LineBuffer1(1583);
--            LineBuffer1(1585) <= LineBuffer1(1584);
--            LineBuffer1(1586) <= LineBuffer1(1585);
--            LineBuffer1(1587) <= LineBuffer1(1586);
--            LineBuffer1(1588) <= LineBuffer1(1587);
--            LineBuffer1(1589) <= LineBuffer1(1588);    
--            LineBuffer1(1590) <= LineBuffer1(1589);
--            LineBuffer1(1591) <= LineBuffer1(1590);
--            LineBuffer1(1592) <= LineBuffer1(1591);
--            LineBuffer1(1593) <= LineBuffer1(1592);
--            LineBuffer1(1594) <= LineBuffer1(1593);
--            LineBuffer1(1595) <= LineBuffer1(1594);
--            LineBuffer1(1596) <= LineBuffer1(1595);
--            LineBuffer1(1597) <= LineBuffer1(1596);
--            LineBuffer1(1598) <= LineBuffer1(1597);
--            LineBuffer1(1599) <= LineBuffer1(1598);    
--            LineBuffer1(1600) <= LineBuffer1(1599);
--            LineBuffer1(1601) <= LineBuffer1(1600);
--            LineBuffer1(1602) <= LineBuffer1(1601);
--            LineBuffer1(1603) <= LineBuffer1(1602);
--            LineBuffer1(1604) <= LineBuffer1(1603);
--            LineBuffer1(1605) <= LineBuffer1(1604);
--            LineBuffer1(1606) <= LineBuffer1(1605);
--            LineBuffer1(1607) <= LineBuffer1(1606);
--            LineBuffer1(1608) <= LineBuffer1(1607);
--            LineBuffer1(1609) <= LineBuffer1(1608);    
--            LineBuffer1(1610) <= LineBuffer1(1609);
--            LineBuffer1(1611) <= LineBuffer1(1610);
--            LineBuffer1(1612) <= LineBuffer1(1611);
--            LineBuffer1(1613) <= LineBuffer1(1612);
--            LineBuffer1(1614) <= LineBuffer1(1613);
--            LineBuffer1(1615) <= LineBuffer1(1614);
--            LineBuffer1(1616) <= LineBuffer1(1615);
--            LineBuffer1(1617) <= LineBuffer1(1616);
--            LineBuffer1(1618) <= LineBuffer1(1617);
--            LineBuffer1(1619) <= LineBuffer1(1618);    
--            LineBuffer1(1620) <= LineBuffer1(1619);
--            LineBuffer1(1621) <= LineBuffer1(1620);
--            LineBuffer1(1622) <= LineBuffer1(1621);
--            LineBuffer1(1623) <= LineBuffer1(1622);
--            LineBuffer1(1624) <= LineBuffer1(1623);
--            LineBuffer1(1625) <= LineBuffer1(1624);
--            LineBuffer1(1626) <= LineBuffer1(1625);
--            LineBuffer1(1627) <= LineBuffer1(1626);
--            LineBuffer1(1628) <= LineBuffer1(1627);
--            LineBuffer1(1629) <= LineBuffer1(1628);    
--            LineBuffer1(1630) <= LineBuffer1(1629);
--            LineBuffer1(1631) <= LineBuffer1(1630);
--            LineBuffer1(1632) <= LineBuffer1(1631);
--            LineBuffer1(1633) <= LineBuffer1(1632);
--            LineBuffer1(1634) <= LineBuffer1(1633);
--            LineBuffer1(1635) <= LineBuffer1(1634);
--            LineBuffer1(1636) <= LineBuffer1(1635);
--            LineBuffer1(1637) <= LineBuffer1(1636);
--            LineBuffer1(1638) <= LineBuffer1(1637);
--            LineBuffer1(1639) <= LineBuffer1(1638);    
--            LineBuffer1(1640) <= LineBuffer1(1639);
--            LineBuffer1(1641) <= LineBuffer1(1640);
--            LineBuffer1(1642) <= LineBuffer1(1641);
--            LineBuffer1(1643) <= LineBuffer1(1642);
--            LineBuffer1(1644) <= LineBuffer1(1643);
--            LineBuffer1(1645) <= LineBuffer1(1644);
--            LineBuffer1(1646) <= LineBuffer1(1645);
--            LineBuffer1(1647) <= LineBuffer1(1646);
--            LineBuffer1(1648) <= LineBuffer1(1647);
--            LineBuffer1(1649) <= LineBuffer1(1648);    
--            LineBuffer1(1650) <= LineBuffer1(1649);
--            LineBuffer1(1651) <= LineBuffer1(1650);
--            LineBuffer1(1652) <= LineBuffer1(1651);
--            LineBuffer1(1653) <= LineBuffer1(1652);
--            LineBuffer1(1654) <= LineBuffer1(1653);
--            LineBuffer1(1655) <= LineBuffer1(1654);
--            LineBuffer1(1656) <= LineBuffer1(1655);
--            LineBuffer1(1657) <= LineBuffer1(1656);
--            LineBuffer1(1658) <= LineBuffer1(1657);
--            LineBuffer1(1659) <= LineBuffer1(1658);    
--            LineBuffer1(1660) <= LineBuffer1(1659);
--            LineBuffer1(1661) <= LineBuffer1(1660);
--            LineBuffer1(1662) <= LineBuffer1(1661);
--            LineBuffer1(1663) <= LineBuffer1(1662);
--            LineBuffer1(1664) <= LineBuffer1(1663);
--            LineBuffer1(1665) <= LineBuffer1(1664);
--            LineBuffer1(1666) <= LineBuffer1(1665);
--            LineBuffer1(1667) <= LineBuffer1(1666);
--            LineBuffer1(1668) <= LineBuffer1(1667);
--            LineBuffer1(1669) <= LineBuffer1(1668);    
--            LineBuffer1(1670) <= LineBuffer1(1669);
--            LineBuffer1(1671) <= LineBuffer1(1670);
--            LineBuffer1(1672) <= LineBuffer1(1671);
--            LineBuffer1(1673) <= LineBuffer1(1672);
--            LineBuffer1(1674) <= LineBuffer1(1673);
--            LineBuffer1(1675) <= LineBuffer1(1674);
--            LineBuffer1(1676) <= LineBuffer1(1675);
--            LineBuffer1(1677) <= LineBuffer1(1676);
--            LineBuffer1(1678) <= LineBuffer1(1677);
--            LineBuffer1(1679) <= LineBuffer1(1678);
--            LineBuffer1(1680) <= LineBuffer1(1679);
--            LineBuffer1(1681) <= LineBuffer1(1680);
--            LineBuffer1(1682) <= LineBuffer1(1681);
--            LineBuffer1(1683) <= LineBuffer1(1682);
--            LineBuffer1(1684) <= LineBuffer1(1683);
--            LineBuffer1(1685) <= LineBuffer1(1684);
--            LineBuffer1(1686) <= LineBuffer1(1685);
--            LineBuffer1(1687) <= LineBuffer1(1686);
--            LineBuffer1(1688) <= LineBuffer1(1687);
--            LineBuffer1(1689) <= LineBuffer1(1688);    
--            LineBuffer1(1690) <= LineBuffer1(1689);
--            LineBuffer1(1691) <= LineBuffer1(1690);
--            LineBuffer1(1692) <= LineBuffer1(1691);
--            LineBuffer1(1693) <= LineBuffer1(1692);
--            LineBuffer1(1694) <= LineBuffer1(1693);
--            LineBuffer1(1695) <= LineBuffer1(1694);
--            LineBuffer1(1696) <= LineBuffer1(1695);
--            LineBuffer1(1697) <= LineBuffer1(1696);
--            LineBuffer1(1698) <= LineBuffer1(1697);
--            LineBuffer1(1699) <= LineBuffer1(1698);    
--            LineBuffer1(1700) <= LineBuffer1(1699);
--            LineBuffer1(1701) <= LineBuffer1(1700);
--            LineBuffer1(1702) <= LineBuffer1(1701);
--            LineBuffer1(1703) <= LineBuffer1(1702);
--            LineBuffer1(1704) <= LineBuffer1(1703);
--            LineBuffer1(1705) <= LineBuffer1(1704);
--            LineBuffer1(1706) <= LineBuffer1(1705);
--            LineBuffer1(1707) <= LineBuffer1(1706);
--            LineBuffer1(1708) <= LineBuffer1(1707);
--            LineBuffer1(1709) <= LineBuffer1(1708);    
--            LineBuffer1(1710) <= LineBuffer1(1709);
--            LineBuffer1(1711) <= LineBuffer1(1710);
--            LineBuffer1(1712) <= LineBuffer1(1711);
--            LineBuffer1(1713) <= LineBuffer1(1712);
--            LineBuffer1(1714) <= LineBuffer1(1713);
--            LineBuffer1(1715) <= LineBuffer1(1714);
--            LineBuffer1(1716) <= LineBuffer1(1715);
--            LineBuffer1(1717) <= LineBuffer1(1716);
--            LineBuffer1(1718) <= LineBuffer1(1717);
--            LineBuffer1(1719) <= LineBuffer1(1718);    
--            LineBuffer1(1720) <= LineBuffer1(1719);
--            LineBuffer1(1721) <= LineBuffer1(1720);
--            LineBuffer1(1722) <= LineBuffer1(1721);
--            LineBuffer1(1723) <= LineBuffer1(1722);
--            LineBuffer1(1724) <= LineBuffer1(1723);
--            LineBuffer1(1725) <= LineBuffer1(1724);
--            LineBuffer1(1726) <= LineBuffer1(1725);
--            LineBuffer1(1727) <= LineBuffer1(1726);
--            LineBuffer1(1728) <= LineBuffer1(1727);
--            LineBuffer1(1729) <= LineBuffer1(1728);    
--            LineBuffer1(1730) <= LineBuffer1(1729);
--            LineBuffer1(1731) <= LineBuffer1(1730);
--            LineBuffer1(1732) <= LineBuffer1(1731);
--            LineBuffer1(1733) <= LineBuffer1(1732);
--            LineBuffer1(1734) <= LineBuffer1(1733);
--            LineBuffer1(1735) <= LineBuffer1(1734);
--            LineBuffer1(1736) <= LineBuffer1(1735);
--            LineBuffer1(1737) <= LineBuffer1(1736);
--            LineBuffer1(1738) <= LineBuffer1(1737);
--            LineBuffer1(1739) <= LineBuffer1(1738);    
--            LineBuffer1(1740) <= LineBuffer1(1739);
--            LineBuffer1(1741) <= LineBuffer1(1740);
--            LineBuffer1(1742) <= LineBuffer1(1741);
--            LineBuffer1(1743) <= LineBuffer1(1742);
--            LineBuffer1(1744) <= LineBuffer1(1743);
--            LineBuffer1(1745) <= LineBuffer1(1744);
--            LineBuffer1(1746) <= LineBuffer1(1745);
--            LineBuffer1(1747) <= LineBuffer1(1746);
--            LineBuffer1(1748) <= LineBuffer1(1747);
--            LineBuffer1(1749) <= LineBuffer1(1748);    
--            LineBuffer1(1750) <= LineBuffer1(1749);
--            LineBuffer1(1751) <= LineBuffer1(1750);
--            LineBuffer1(1752) <= LineBuffer1(1751);
--            LineBuffer1(1753) <= LineBuffer1(1752);
--            LineBuffer1(1754) <= LineBuffer1(1753);
--            LineBuffer1(1755) <= LineBuffer1(1754);
--            LineBuffer1(1756) <= LineBuffer1(1755);
--            LineBuffer1(1757) <= LineBuffer1(1756);
--            LineBuffer1(1758) <= LineBuffer1(1757);
--            LineBuffer1(1759) <= LineBuffer1(1758);    
--            LineBuffer1(1760) <= LineBuffer1(1759);
--            LineBuffer1(1761) <= LineBuffer1(1760);
--            LineBuffer1(1762) <= LineBuffer1(1761);
--            LineBuffer1(1763) <= LineBuffer1(1762);
--            LineBuffer1(1764) <= LineBuffer1(1763);
--            LineBuffer1(1765) <= LineBuffer1(1764);
--            LineBuffer1(1766) <= LineBuffer1(1765);
--            LineBuffer1(1767) <= LineBuffer1(1766);
--            LineBuffer1(1768) <= LineBuffer1(1767);
--            LineBuffer1(1769) <= LineBuffer1(1768);    
--            LineBuffer1(1770) <= LineBuffer1(1769);
--            LineBuffer1(1771) <= LineBuffer1(1770);
--            LineBuffer1(1772) <= LineBuffer1(1771);
--            LineBuffer1(1773) <= LineBuffer1(1772);
--            LineBuffer1(1774) <= LineBuffer1(1773);
--            LineBuffer1(1775) <= LineBuffer1(1774);
--            LineBuffer1(1776) <= LineBuffer1(1775);
--            LineBuffer1(1777) <= LineBuffer1(1776);
--            LineBuffer1(1778) <= LineBuffer1(1777);
--            LineBuffer1(1779) <= LineBuffer1(1778);
--            LineBuffer1(1780) <= LineBuffer1(1779);
--            LineBuffer1(1781) <= LineBuffer1(1780);
--            LineBuffer1(1782) <= LineBuffer1(1781);
--            LineBuffer1(1783) <= LineBuffer1(1782);
--            LineBuffer1(1784) <= LineBuffer1(1783);
--            LineBuffer1(1785) <= LineBuffer1(1784);
--            LineBuffer1(1786) <= LineBuffer1(1785);
--            LineBuffer1(1787) <= LineBuffer1(1786);
--            LineBuffer1(1788) <= LineBuffer1(1787);
--            LineBuffer1(1789) <= LineBuffer1(1788);    
--            LineBuffer1(1790) <= LineBuffer1(1789);
--            LineBuffer1(1791) <= LineBuffer1(1790);
--            LineBuffer1(1792) <= LineBuffer1(1791);
--            LineBuffer1(1793) <= LineBuffer1(1792);
--            LineBuffer1(1794) <= LineBuffer1(1793);
--            LineBuffer1(1795) <= LineBuffer1(1794);
--            LineBuffer1(1796) <= LineBuffer1(1795);
--            LineBuffer1(1797) <= LineBuffer1(1796);
--            LineBuffer1(1798) <= LineBuffer1(1797);
--            LineBuffer1(1799) <= LineBuffer1(1798);    
--            LineBuffer1(1800) <= LineBuffer1(1799);
--            LineBuffer1(1801) <= LineBuffer1(1800);
--            LineBuffer1(1802) <= LineBuffer1(1801);
--            LineBuffer1(1803) <= LineBuffer1(1802);
--            LineBuffer1(1804) <= LineBuffer1(1803);
--            LineBuffer1(1805) <= LineBuffer1(1804);
--            LineBuffer1(1806) <= LineBuffer1(1805);
--            LineBuffer1(1807) <= LineBuffer1(1806);
--            LineBuffer1(1808) <= LineBuffer1(1807);
--            LineBuffer1(1809) <= LineBuffer1(1808);    
--            LineBuffer1(1810) <= LineBuffer1(1809);
--            LineBuffer1(1811) <= LineBuffer1(1810);
--            LineBuffer1(1812) <= LineBuffer1(1811);
--            LineBuffer1(1813) <= LineBuffer1(1812);
--            LineBuffer1(1814) <= LineBuffer1(1813);
--            LineBuffer1(1815) <= LineBuffer1(1814);
--            LineBuffer1(1816) <= LineBuffer1(1815);
--            LineBuffer1(1817) <= LineBuffer1(1816);
--            LineBuffer1(1818) <= LineBuffer1(1817);
--            LineBuffer1(1819) <= LineBuffer1(1818);    
--            LineBuffer1(1820) <= LineBuffer1(1819);
--            LineBuffer1(1821) <= LineBuffer1(1820);
--            LineBuffer1(1822) <= LineBuffer1(1821);
--            LineBuffer1(1823) <= LineBuffer1(1822);
--            LineBuffer1(1824) <= LineBuffer1(1823);
--            LineBuffer1(1825) <= LineBuffer1(1824);
--            LineBuffer1(1826) <= LineBuffer1(1825);
--            LineBuffer1(1827) <= LineBuffer1(1826);
--            LineBuffer1(1828) <= LineBuffer1(1827);
--            LineBuffer1(1829) <= LineBuffer1(1828);    
--            LineBuffer1(1830) <= LineBuffer1(1829);
--            LineBuffer1(1831) <= LineBuffer1(1830);
--            LineBuffer1(1832) <= LineBuffer1(1831);
--            LineBuffer1(1833) <= LineBuffer1(1832);
--            LineBuffer1(1834) <= LineBuffer1(1833);
--            LineBuffer1(1835) <= LineBuffer1(1834);
--            LineBuffer1(1836) <= LineBuffer1(1835);
--            LineBuffer1(1837) <= LineBuffer1(1836);
--            LineBuffer1(1838) <= LineBuffer1(1837);
--            LineBuffer1(1839) <= LineBuffer1(1838);    
--            LineBuffer1(1840) <= LineBuffer1(1839);
--            LineBuffer1(1841) <= LineBuffer1(1840);
--            LineBuffer1(1842) <= LineBuffer1(1841);
--            LineBuffer1(1843) <= LineBuffer1(1842);
--            LineBuffer1(1844) <= LineBuffer1(1843);
--            LineBuffer1(1845) <= LineBuffer1(1844);
--            LineBuffer1(1846) <= LineBuffer1(1845);
--            LineBuffer1(1847) <= LineBuffer1(1846);
--            LineBuffer1(1848) <= LineBuffer1(1847);
--            LineBuffer1(1849) <= LineBuffer1(1848);    
--            LineBuffer1(1850) <= LineBuffer1(1849);
--            LineBuffer1(1851) <= LineBuffer1(1850);
--            LineBuffer1(1852) <= LineBuffer1(1851);
--            LineBuffer1(1853) <= LineBuffer1(1852);
--            LineBuffer1(1854) <= LineBuffer1(1853);
--            LineBuffer1(1855) <= LineBuffer1(1854);
--            LineBuffer1(1856) <= LineBuffer1(1855);
--            LineBuffer1(1857) <= LineBuffer1(1856);
--            LineBuffer1(1858) <= LineBuffer1(1857);
--            LineBuffer1(1859) <= LineBuffer1(1858);    
--            LineBuffer1(1860) <= LineBuffer1(1859);
--            LineBuffer1(1861) <= LineBuffer1(1860);
--            LineBuffer1(1862) <= LineBuffer1(1861);
--            LineBuffer1(1863) <= LineBuffer1(1862);
--            LineBuffer1(1864) <= LineBuffer1(1863);
--            LineBuffer1(1865) <= LineBuffer1(1864);
--            LineBuffer1(1866) <= LineBuffer1(1865);
--            LineBuffer1(1867) <= LineBuffer1(1866);
--            LineBuffer1(1868) <= LineBuffer1(1867);
--            LineBuffer1(1869) <= LineBuffer1(1868);    
--            LineBuffer1(1870) <= LineBuffer1(1869);
--            LineBuffer1(1871) <= LineBuffer1(1870);
--            LineBuffer1(1872) <= LineBuffer1(1871);
--            LineBuffer1(1873) <= LineBuffer1(1872);
--            LineBuffer1(1874) <= LineBuffer1(1873);
--            LineBuffer1(1875) <= LineBuffer1(1874);
--            LineBuffer1(1876) <= LineBuffer1(1875);
--            LineBuffer1(1877) <= LineBuffer1(1876);
--            LineBuffer1(1878) <= LineBuffer1(1877);
--            LineBuffer1(1879) <= LineBuffer1(1878);
--            LineBuffer1(1880) <= LineBuffer1(1879);
--            LineBuffer1(1881) <= LineBuffer1(1880);
--            LineBuffer1(1882) <= LineBuffer1(1881);
--            LineBuffer1(1883) <= LineBuffer1(1882);
--            LineBuffer1(1884) <= LineBuffer1(1883);
--            LineBuffer1(1885) <= LineBuffer1(1884);
--            LineBuffer1(1886) <= LineBuffer1(1885);
--            LineBuffer1(1887) <= LineBuffer1(1886);
--            LineBuffer1(1888) <= LineBuffer1(1887);
--            LineBuffer1(1889) <= LineBuffer1(1888);    
--            LineBuffer1(1890) <= LineBuffer1(1889);
--            LineBuffer1(1891) <= LineBuffer1(1890);
--            LineBuffer1(1892) <= LineBuffer1(1891);
--            LineBuffer1(1893) <= LineBuffer1(1892);
--            LineBuffer1(1894) <= LineBuffer1(1893);
--            LineBuffer1(1895) <= LineBuffer1(1894);
--            LineBuffer1(1896) <= LineBuffer1(1895);
--            LineBuffer1(1897) <= LineBuffer1(1896);
--            LineBuffer1(1898) <= LineBuffer1(1897);
--            LineBuffer1(1899) <= LineBuffer1(1898);    
--            LineBuffer1(1900) <= LineBuffer1(1899);
--            LineBuffer1(1901) <= LineBuffer1(1900);
--            LineBuffer1(1902) <= LineBuffer1(1901);
--            LineBuffer1(1903) <= LineBuffer1(1902);
--            LineBuffer1(1904) <= LineBuffer1(1903);
--            LineBuffer1(1905) <= LineBuffer1(1904);
--            LineBuffer1(1906) <= LineBuffer1(1905);
--            LineBuffer1(1907) <= LineBuffer1(1906);
--            LineBuffer1(1908) <= LineBuffer1(1907);
--            LineBuffer1(1909) <= LineBuffer1(1908);    
--            LineBuffer1(1910) <= LineBuffer1(1909);
--            LineBuffer1(1911) <= LineBuffer1(1910);
--            LineBuffer1(1912) <= LineBuffer1(1911);
--            LineBuffer1(1913) <= LineBuffer1(1912);
--            LineBuffer1(1914) <= LineBuffer1(1913);
--            LineBuffer1(1915) <= LineBuffer1(1914);
--            LineBuffer1(1916) <= LineBuffer1(1915);
--            LineBuffer1(1917) <= LineBuffer1(1916);
--            LineBuffer1(1918) <= LineBuffer1(1917);
--            LineBuffer1(1919) <= LineBuffer1(1918);	

			
			
			
			LineBuffer2(0) <= LineBuffer1(1279);
			LineBuffer2(1) <= LineBuffer2(0);
			LineBuffer2(2) <= LineBuffer2(1);
			LineBuffer2(3) <= LineBuffer2(2);
			LineBuffer2(4) <= LineBuffer2(3);
			LineBuffer2(5) <= LineBuffer2(4);
			LineBuffer2(6) <= LineBuffer2(5);
			LineBuffer2(7) <= LineBuffer2(6);
			LineBuffer2(8) <= LineBuffer2(7);
			LineBuffer2(9) <= LineBuffer2(8);	
			LineBuffer2(10) <= LineBuffer2(9);
			LineBuffer2(11) <= LineBuffer2(10);
			LineBuffer2(12) <= LineBuffer2(11);
			LineBuffer2(13) <= LineBuffer2(12);
			LineBuffer2(14) <= LineBuffer2(13);
			LineBuffer2(15) <= LineBuffer2(14);
			LineBuffer2(16) <= LineBuffer2(15);
			LineBuffer2(17) <= LineBuffer2(16);
			LineBuffer2(18) <= LineBuffer2(17);
			LineBuffer2(19) <= LineBuffer2(18);	
			LineBuffer2(20) <= LineBuffer2(19);
			LineBuffer2(21) <= LineBuffer2(20);
			LineBuffer2(22) <= LineBuffer2(21);
			LineBuffer2(23) <= LineBuffer2(22);
			LineBuffer2(24) <= LineBuffer2(23);
			LineBuffer2(25) <= LineBuffer2(24);
			LineBuffer2(26) <= LineBuffer2(25);
			LineBuffer2(27) <= LineBuffer2(26);
			LineBuffer2(28) <= LineBuffer2(27);
			LineBuffer2(29) <= LineBuffer2(28);	
			LineBuffer2(30) <= LineBuffer2(29);
			LineBuffer2(31) <= LineBuffer2(30);
			LineBuffer2(32) <= LineBuffer2(31);
			LineBuffer2(33) <= LineBuffer2(32);
			LineBuffer2(34) <= LineBuffer2(33);
			LineBuffer2(35) <= LineBuffer2(34);
			LineBuffer2(36) <= LineBuffer2(35);
			LineBuffer2(37) <= LineBuffer2(36);
			LineBuffer2(38) <= LineBuffer2(37);
			LineBuffer2(39) <= LineBuffer2(38);	
			LineBuffer2(40) <= LineBuffer2(39);
			LineBuffer2(41) <= LineBuffer2(40);
			LineBuffer2(42) <= LineBuffer2(41);
			LineBuffer2(43) <= LineBuffer2(42);
			LineBuffer2(44) <= LineBuffer2(43);
			LineBuffer2(45) <= LineBuffer2(44);
			LineBuffer2(46) <= LineBuffer2(45);
			LineBuffer2(47) <= LineBuffer2(46);
			LineBuffer2(48) <= LineBuffer2(47);
			LineBuffer2(49) <= LineBuffer2(48);	
			LineBuffer2(50) <= LineBuffer2(49);
			LineBuffer2(51) <= LineBuffer2(50);
			LineBuffer2(52) <= LineBuffer2(51);
			LineBuffer2(53) <= LineBuffer2(52);
			LineBuffer2(54) <= LineBuffer2(53);
			LineBuffer2(55) <= LineBuffer2(54);
			LineBuffer2(56) <= LineBuffer2(55);
			LineBuffer2(57) <= LineBuffer2(56);
			LineBuffer2(58) <= LineBuffer2(57);
			LineBuffer2(59) <= LineBuffer2(58);	
			LineBuffer2(60) <= LineBuffer2(59);
			LineBuffer2(61) <= LineBuffer2(60);
			LineBuffer2(62) <= LineBuffer2(61);
			LineBuffer2(63) <= LineBuffer2(62);
			LineBuffer2(64) <= LineBuffer2(63);
			LineBuffer2(65) <= LineBuffer2(64);
			LineBuffer2(66) <= LineBuffer2(65);
			LineBuffer2(67) <= LineBuffer2(66);
			LineBuffer2(68) <= LineBuffer2(67);
			LineBuffer2(69) <= LineBuffer2(68);	
			LineBuffer2(70) <= LineBuffer2(69);
			LineBuffer2(71) <= LineBuffer2(70);
			LineBuffer2(72) <= LineBuffer2(71);
			LineBuffer2(73) <= LineBuffer2(72);
			LineBuffer2(74) <= LineBuffer2(73);
			LineBuffer2(75) <= LineBuffer2(74);
			LineBuffer2(76) <= LineBuffer2(75);
			LineBuffer2(77) <= LineBuffer2(76);
			LineBuffer2(78) <= LineBuffer2(77);
			LineBuffer2(79) <= LineBuffer2(78);	
			LineBuffer2(80) <= LineBuffer2(79);
			LineBuffer2(81) <= LineBuffer2(80);
			LineBuffer2(82) <= LineBuffer2(81);
			LineBuffer2(83) <= LineBuffer2(82);
			LineBuffer2(84) <= LineBuffer2(83);
			LineBuffer2(85) <= LineBuffer2(84);
			LineBuffer2(86) <= LineBuffer2(85);
			LineBuffer2(87) <= LineBuffer2(86);
			LineBuffer2(88) <= LineBuffer2(87);
			LineBuffer2(89) <= LineBuffer2(88);	
			LineBuffer2(90) <= LineBuffer2(89);
			LineBuffer2(91) <= LineBuffer2(90);
			LineBuffer2(92) <= LineBuffer2(91);
			LineBuffer2(93) <= LineBuffer2(92);
			LineBuffer2(94) <= LineBuffer2(93);
			LineBuffer2(95) <= LineBuffer2(94);
			LineBuffer2(96) <= LineBuffer2(95);
			LineBuffer2(97) <= LineBuffer2(96);
			LineBuffer2(98) <= LineBuffer2(97);
			LineBuffer2(99) <= LineBuffer2(98);	
			LineBuffer2(100) <= LineBuffer2(99);
			LineBuffer2(101) <= LineBuffer2(100);
			LineBuffer2(102) <= LineBuffer2(101);
			LineBuffer2(103) <= LineBuffer2(102);
			LineBuffer2(104) <= LineBuffer2(103);
			LineBuffer2(105) <= LineBuffer2(104);
			LineBuffer2(106) <= LineBuffer2(105);
			LineBuffer2(107) <= LineBuffer2(106);
			LineBuffer2(108) <= LineBuffer2(107);
			LineBuffer2(109) <= LineBuffer2(108);	
			LineBuffer2(110) <= LineBuffer2(109);
			LineBuffer2(111) <= LineBuffer2(110);
			LineBuffer2(112) <= LineBuffer2(111);
			LineBuffer2(113) <= LineBuffer2(112);
			LineBuffer2(114) <= LineBuffer2(113);
			LineBuffer2(115) <= LineBuffer2(114);
			LineBuffer2(116) <= LineBuffer2(115);
			LineBuffer2(117) <= LineBuffer2(116);
			LineBuffer2(118) <= LineBuffer2(117);
			LineBuffer2(119) <= LineBuffer2(118);	
			LineBuffer2(120) <= LineBuffer2(119);
			LineBuffer2(121) <= LineBuffer2(120);
			LineBuffer2(122) <= LineBuffer2(121);
			LineBuffer2(123) <= LineBuffer2(122);
			LineBuffer2(124) <= LineBuffer2(123);
			LineBuffer2(125) <= LineBuffer2(124);
			LineBuffer2(126) <= LineBuffer2(125);
			LineBuffer2(127) <= LineBuffer2(126);
			LineBuffer2(128) <= LineBuffer2(127);
			LineBuffer2(129) <= LineBuffer2(128);	
			LineBuffer2(130) <= LineBuffer2(129);
			LineBuffer2(131) <= LineBuffer2(130);
			LineBuffer2(132) <= LineBuffer2(131);
			LineBuffer2(133) <= LineBuffer2(132);
			LineBuffer2(134) <= LineBuffer2(133);
			LineBuffer2(135) <= LineBuffer2(134);
			LineBuffer2(136) <= LineBuffer2(135);
			LineBuffer2(137) <= LineBuffer2(136);
			LineBuffer2(138) <= LineBuffer2(137);
			LineBuffer2(139) <= LineBuffer2(138);	
			LineBuffer2(140) <= LineBuffer2(139);
			LineBuffer2(141) <= LineBuffer2(140);
			LineBuffer2(142) <= LineBuffer2(141);
			LineBuffer2(143) <= LineBuffer2(142);
			LineBuffer2(144) <= LineBuffer2(143);
			LineBuffer2(145) <= LineBuffer2(144);
			LineBuffer2(146) <= LineBuffer2(145);
			LineBuffer2(147) <= LineBuffer2(146);
			LineBuffer2(148) <= LineBuffer2(147);
			LineBuffer2(149) <= LineBuffer2(148);	
			LineBuffer2(150) <= LineBuffer2(149);
			LineBuffer2(151) <= LineBuffer2(150);
			LineBuffer2(152) <= LineBuffer2(151);
			LineBuffer2(153) <= LineBuffer2(152);
			LineBuffer2(154) <= LineBuffer2(153);
			LineBuffer2(155) <= LineBuffer2(154);
			LineBuffer2(156) <= LineBuffer2(155);
			LineBuffer2(157) <= LineBuffer2(156);
			LineBuffer2(158) <= LineBuffer2(157);
			LineBuffer2(159) <= LineBuffer2(158);	
			LineBuffer2(160) <= LineBuffer2(159);
			LineBuffer2(161) <= LineBuffer2(160);
			LineBuffer2(162) <= LineBuffer2(161);
			LineBuffer2(163) <= LineBuffer2(162);
			LineBuffer2(164) <= LineBuffer2(163);
			LineBuffer2(165) <= LineBuffer2(164);
			LineBuffer2(166) <= LineBuffer2(165);
			LineBuffer2(167) <= LineBuffer2(166);
			LineBuffer2(168) <= LineBuffer2(167);
			LineBuffer2(169) <= LineBuffer2(168);	
			LineBuffer2(170) <= LineBuffer2(169);
			LineBuffer2(171) <= LineBuffer2(170);
			LineBuffer2(172) <= LineBuffer2(171);
			LineBuffer2(173) <= LineBuffer2(172);
			LineBuffer2(174) <= LineBuffer2(173);
			LineBuffer2(175) <= LineBuffer2(174);
			LineBuffer2(176) <= LineBuffer2(175);
			LineBuffer2(177) <= LineBuffer2(176);
			LineBuffer2(178) <= LineBuffer2(177);
			LineBuffer2(179) <= LineBuffer2(178);	
			LineBuffer2(180) <= LineBuffer2(179);
			LineBuffer2(181) <= LineBuffer2(180);
			LineBuffer2(182) <= LineBuffer2(181);
			LineBuffer2(183) <= LineBuffer2(182);
			LineBuffer2(184) <= LineBuffer2(183);
			LineBuffer2(185) <= LineBuffer2(184);
			LineBuffer2(186) <= LineBuffer2(185);
			LineBuffer2(187) <= LineBuffer2(186);
			LineBuffer2(188) <= LineBuffer2(187);
			LineBuffer2(189) <= LineBuffer2(188);	
			LineBuffer2(190) <= LineBuffer2(189);
			LineBuffer2(191) <= LineBuffer2(190);
			LineBuffer2(192) <= LineBuffer2(191);
			LineBuffer2(193) <= LineBuffer2(192);
			LineBuffer2(194) <= LineBuffer2(193);
			LineBuffer2(195) <= LineBuffer2(194);
			LineBuffer2(196) <= LineBuffer2(195);
			LineBuffer2(197) <= LineBuffer2(196);
			LineBuffer2(198) <= LineBuffer2(197);
			LineBuffer2(199) <= LineBuffer2(198);
			LineBuffer2(200) <= LineBuffer2(199);
			LineBuffer2(201) <= LineBuffer2(200);
			LineBuffer2(202) <= LineBuffer2(201);
			LineBuffer2(203) <= LineBuffer2(202);
			LineBuffer2(204) <= LineBuffer2(203);
			LineBuffer2(205) <= LineBuffer2(204);
			LineBuffer2(206) <= LineBuffer2(205);
			LineBuffer2(207) <= LineBuffer2(206);
			LineBuffer2(208) <= LineBuffer2(207);
			LineBuffer2(209) <= LineBuffer2(208);	
			LineBuffer2(210) <= LineBuffer2(209);
			LineBuffer2(211) <= LineBuffer2(210);
			LineBuffer2(212) <= LineBuffer2(211);
			LineBuffer2(213) <= LineBuffer2(212);
			LineBuffer2(214) <= LineBuffer2(213);
			LineBuffer2(215) <= LineBuffer2(214);
			LineBuffer2(216) <= LineBuffer2(215);
			LineBuffer2(217) <= LineBuffer2(216);
			LineBuffer2(218) <= LineBuffer2(217);
			LineBuffer2(219) <= LineBuffer2(218);	
			LineBuffer2(220) <= LineBuffer2(219);
			LineBuffer2(221) <= LineBuffer2(220);
			LineBuffer2(222) <= LineBuffer2(221);
			LineBuffer2(223) <= LineBuffer2(222);
			LineBuffer2(224) <= LineBuffer2(223);
			LineBuffer2(225) <= LineBuffer2(224);
			LineBuffer2(226) <= LineBuffer2(225);
			LineBuffer2(227) <= LineBuffer2(226);
			LineBuffer2(228) <= LineBuffer2(227);
			LineBuffer2(229) <= LineBuffer2(228);	
			LineBuffer2(230) <= LineBuffer2(229);
			LineBuffer2(231) <= LineBuffer2(230);
			LineBuffer2(232) <= LineBuffer2(231);
			LineBuffer2(233) <= LineBuffer2(232);
			LineBuffer2(234) <= LineBuffer2(233);
			LineBuffer2(235) <= LineBuffer2(234);
			LineBuffer2(236) <= LineBuffer2(235);
			LineBuffer2(237) <= LineBuffer2(236);
			LineBuffer2(238) <= LineBuffer2(237);
			LineBuffer2(239) <= LineBuffer2(238);	
			LineBuffer2(240) <= LineBuffer2(239);
			LineBuffer2(241) <= LineBuffer2(240);
			LineBuffer2(242) <= LineBuffer2(241);
			LineBuffer2(243) <= LineBuffer2(242);
			LineBuffer2(244) <= LineBuffer2(243);
			LineBuffer2(245) <= LineBuffer2(244);
			LineBuffer2(246) <= LineBuffer2(245);
			LineBuffer2(247) <= LineBuffer2(246);
			LineBuffer2(248) <= LineBuffer2(247);
			LineBuffer2(249) <= LineBuffer2(248);	
			LineBuffer2(250) <= LineBuffer2(249);
			LineBuffer2(251) <= LineBuffer2(250);
			LineBuffer2(252) <= LineBuffer2(251);
			LineBuffer2(253) <= LineBuffer2(252);
			LineBuffer2(254) <= LineBuffer2(253);
			LineBuffer2(255) <= LineBuffer2(254);
			LineBuffer2(256) <= LineBuffer2(255);
			LineBuffer2(257) <= LineBuffer2(256);
			LineBuffer2(258) <= LineBuffer2(257);
			LineBuffer2(259) <= LineBuffer2(258);	
			LineBuffer2(260) <= LineBuffer2(259);
			LineBuffer2(261) <= LineBuffer2(260);
			LineBuffer2(262) <= LineBuffer2(261);
			LineBuffer2(263) <= LineBuffer2(262);
			LineBuffer2(264) <= LineBuffer2(263);
			LineBuffer2(265) <= LineBuffer2(264);
			LineBuffer2(266) <= LineBuffer2(265);
			LineBuffer2(267) <= LineBuffer2(266);
			LineBuffer2(268) <= LineBuffer2(267);
			LineBuffer2(269) <= LineBuffer2(268);	
			LineBuffer2(270) <= LineBuffer2(269);
			LineBuffer2(271) <= LineBuffer2(270);
			LineBuffer2(272) <= LineBuffer2(271);
			LineBuffer2(273) <= LineBuffer2(272);
			LineBuffer2(274) <= LineBuffer2(273);
			LineBuffer2(275) <= LineBuffer2(274);
			LineBuffer2(276) <= LineBuffer2(275);
			LineBuffer2(277) <= LineBuffer2(276);
			LineBuffer2(278) <= LineBuffer2(277);
			LineBuffer2(279) <= LineBuffer2(278);	
			LineBuffer2(280) <= LineBuffer2(279);
			LineBuffer2(281) <= LineBuffer2(280);
			LineBuffer2(282) <= LineBuffer2(281);
			LineBuffer2(283) <= LineBuffer2(282);
			LineBuffer2(284) <= LineBuffer2(283);
			LineBuffer2(285) <= LineBuffer2(284);
			LineBuffer2(286) <= LineBuffer2(285);
			LineBuffer2(287) <= LineBuffer2(286);
			LineBuffer2(288) <= LineBuffer2(287);
			LineBuffer2(289) <= LineBuffer2(288);	
			LineBuffer2(290) <= LineBuffer2(289);
			LineBuffer2(291) <= LineBuffer2(290);
			LineBuffer2(292) <= LineBuffer2(291);
			LineBuffer2(293) <= LineBuffer2(292);
			LineBuffer2(294) <= LineBuffer2(293);
			LineBuffer2(295) <= LineBuffer2(294);
			LineBuffer2(296) <= LineBuffer2(295);
			LineBuffer2(297) <= LineBuffer2(296);
			LineBuffer2(298) <= LineBuffer2(297);
			LineBuffer2(299) <= LineBuffer2(298);	
			LineBuffer2(300) <= LineBuffer2(299);	
			LineBuffer2(301) <= LineBuffer2(300);
			LineBuffer2(302) <= LineBuffer2(301);
			LineBuffer2(303) <= LineBuffer2(302);
			LineBuffer2(304) <= LineBuffer2(303);
			LineBuffer2(305) <= LineBuffer2(304);
			LineBuffer2(306) <= LineBuffer2(305);
			LineBuffer2(307) <= LineBuffer2(306);
			LineBuffer2(308) <= LineBuffer2(307);
			LineBuffer2(309) <= LineBuffer2(308);	
			LineBuffer2(310) <= LineBuffer2(309);
			LineBuffer2(311) <= LineBuffer2(310);
			LineBuffer2(312) <= LineBuffer2(311);
			LineBuffer2(313) <= LineBuffer2(312);
			LineBuffer2(314) <= LineBuffer2(313);
			LineBuffer2(315) <= LineBuffer2(314);
			LineBuffer2(316) <= LineBuffer2(315);
			LineBuffer2(317) <= LineBuffer2(316);
			LineBuffer2(318) <= LineBuffer2(317);
			LineBuffer2(319) <= LineBuffer2(318);	
			LineBuffer2(320) <= LineBuffer2(319);
			LineBuffer2(321) <= LineBuffer2(320);
			LineBuffer2(322) <= LineBuffer2(321);
			LineBuffer2(323) <= LineBuffer2(322);
			LineBuffer2(324) <= LineBuffer2(323);
			LineBuffer2(325) <= LineBuffer2(324);
			LineBuffer2(326) <= LineBuffer2(325);
			LineBuffer2(327) <= LineBuffer2(326);
			LineBuffer2(328) <= LineBuffer2(327);
			LineBuffer2(329) <= LineBuffer2(328);	
			LineBuffer2(330) <= LineBuffer2(329);
			LineBuffer2(331) <= LineBuffer2(330);
			LineBuffer2(332) <= LineBuffer2(331);
			LineBuffer2(333) <= LineBuffer2(332);
			LineBuffer2(334) <= LineBuffer2(333);
			LineBuffer2(335) <= LineBuffer2(334);
			LineBuffer2(336) <= LineBuffer2(335);
			LineBuffer2(337) <= LineBuffer2(336);
			LineBuffer2(338) <= LineBuffer2(337);
			LineBuffer2(339) <= LineBuffer2(338);	
			LineBuffer2(340) <= LineBuffer2(339);
			LineBuffer2(341) <= LineBuffer2(340);
			LineBuffer2(342) <= LineBuffer2(341);
			LineBuffer2(343) <= LineBuffer2(342);
			LineBuffer2(344) <= LineBuffer2(343);
			LineBuffer2(345) <= LineBuffer2(344);
			LineBuffer2(346) <= LineBuffer2(345);
			LineBuffer2(347) <= LineBuffer2(346);
			LineBuffer2(348) <= LineBuffer2(347);
			LineBuffer2(349) <= LineBuffer2(348);	
			LineBuffer2(350) <= LineBuffer2(349);
			LineBuffer2(351) <= LineBuffer2(350);
			LineBuffer2(352) <= LineBuffer2(351);
			LineBuffer2(353) <= LineBuffer2(352);
			LineBuffer2(354) <= LineBuffer2(353);
			LineBuffer2(355) <= LineBuffer2(354);
			LineBuffer2(356) <= LineBuffer2(355);
			LineBuffer2(357) <= LineBuffer2(356);
			LineBuffer2(358) <= LineBuffer2(357);
			LineBuffer2(359) <= LineBuffer2(358);	
			LineBuffer2(360) <= LineBuffer2(359);
			LineBuffer2(361) <= LineBuffer2(360);
			LineBuffer2(362) <= LineBuffer2(361);
			LineBuffer2(363) <= LineBuffer2(362);
			LineBuffer2(364) <= LineBuffer2(363);
			LineBuffer2(365) <= LineBuffer2(364);
			LineBuffer2(366) <= LineBuffer2(365);
			LineBuffer2(367) <= LineBuffer2(366);
			LineBuffer2(368) <= LineBuffer2(367);
			LineBuffer2(369) <= LineBuffer2(368);	
			LineBuffer2(370) <= LineBuffer2(369);
			LineBuffer2(371) <= LineBuffer2(370);
			LineBuffer2(372) <= LineBuffer2(371);
			LineBuffer2(373) <= LineBuffer2(372);
			LineBuffer2(374) <= LineBuffer2(373);
			LineBuffer2(375) <= LineBuffer2(374);
			LineBuffer2(376) <= LineBuffer2(375);
			LineBuffer2(377) <= LineBuffer2(376);
			LineBuffer2(378) <= LineBuffer2(377);
			LineBuffer2(379) <= LineBuffer2(378);	
			LineBuffer2(380) <= LineBuffer2(379);
			LineBuffer2(381) <= LineBuffer2(380);
			LineBuffer2(382) <= LineBuffer2(381);
			LineBuffer2(383) <= LineBuffer2(382);
			LineBuffer2(384) <= LineBuffer2(383);
			LineBuffer2(385) <= LineBuffer2(384);
			LineBuffer2(386) <= LineBuffer2(385);
			LineBuffer2(387) <= LineBuffer2(386);
			LineBuffer2(388) <= LineBuffer2(387);
			LineBuffer2(389) <= LineBuffer2(388);	
			LineBuffer2(390) <= LineBuffer2(389);
			LineBuffer2(391) <= LineBuffer2(390);
			LineBuffer2(392) <= LineBuffer2(391);
			LineBuffer2(393) <= LineBuffer2(392);
			LineBuffer2(394) <= LineBuffer2(393);
			LineBuffer2(395) <= LineBuffer2(394);
			LineBuffer2(396) <= LineBuffer2(395);
			LineBuffer2(397) <= LineBuffer2(396);
			LineBuffer2(398) <= LineBuffer2(397);
			LineBuffer2(399) <= LineBuffer2(398);
			LineBuffer2(400) <= LineBuffer2(399);	
			LineBuffer2(401) <= LineBuffer2(400);
			LineBuffer2(402) <= LineBuffer2(401);
			LineBuffer2(403) <= LineBuffer2(402);
			LineBuffer2(404) <= LineBuffer2(403);
			LineBuffer2(405) <= LineBuffer2(404);
			LineBuffer2(406) <= LineBuffer2(405);
			LineBuffer2(407) <= LineBuffer2(406);
			LineBuffer2(408) <= LineBuffer2(407);
			LineBuffer2(409) <= LineBuffer2(408);	
			LineBuffer2(410) <= LineBuffer2(409);
			LineBuffer2(411) <= LineBuffer2(410);
			LineBuffer2(412) <= LineBuffer2(411);
			LineBuffer2(413) <= LineBuffer2(412);
			LineBuffer2(414) <= LineBuffer2(413);
			LineBuffer2(415) <= LineBuffer2(414);
			LineBuffer2(416) <= LineBuffer2(415);
			LineBuffer2(417) <= LineBuffer2(416);
			LineBuffer2(418) <= LineBuffer2(417);
			LineBuffer2(419) <= LineBuffer2(418);	
			LineBuffer2(420) <= LineBuffer2(419);
			LineBuffer2(421) <= LineBuffer2(420);
			LineBuffer2(422) <= LineBuffer2(421);
			LineBuffer2(423) <= LineBuffer2(422);
			LineBuffer2(424) <= LineBuffer2(423);
			LineBuffer2(425) <= LineBuffer2(424);
			LineBuffer2(426) <= LineBuffer2(425);
			LineBuffer2(427) <= LineBuffer2(426);
			LineBuffer2(428) <= LineBuffer2(427);
			LineBuffer2(429) <= LineBuffer2(428);	
			LineBuffer2(430) <= LineBuffer2(429);
			LineBuffer2(431) <= LineBuffer2(430);
			LineBuffer2(432) <= LineBuffer2(431);
			LineBuffer2(433) <= LineBuffer2(432);
			LineBuffer2(434) <= LineBuffer2(433);
			LineBuffer2(435) <= LineBuffer2(434);
			LineBuffer2(436) <= LineBuffer2(435);
			LineBuffer2(437) <= LineBuffer2(436);
			LineBuffer2(438) <= LineBuffer2(437);
			LineBuffer2(439) <= LineBuffer2(438);	
			LineBuffer2(440) <= LineBuffer2(439);
			LineBuffer2(441) <= LineBuffer2(440);
			LineBuffer2(442) <= LineBuffer2(441);
			LineBuffer2(443) <= LineBuffer2(442);
			LineBuffer2(444) <= LineBuffer2(443);
			LineBuffer2(445) <= LineBuffer2(444);
			LineBuffer2(446) <= LineBuffer2(445);
			LineBuffer2(447) <= LineBuffer2(446);
			LineBuffer2(448) <= LineBuffer2(447);
			LineBuffer2(449) <= LineBuffer2(448);	
			LineBuffer2(450) <= LineBuffer2(449);
			LineBuffer2(451) <= LineBuffer2(450);
			LineBuffer2(452) <= LineBuffer2(451);
			LineBuffer2(453) <= LineBuffer2(452);
			LineBuffer2(454) <= LineBuffer2(453);
			LineBuffer2(455) <= LineBuffer2(454);
			LineBuffer2(456) <= LineBuffer2(455);
			LineBuffer2(457) <= LineBuffer2(456);
			LineBuffer2(458) <= LineBuffer2(457);
			LineBuffer2(459) <= LineBuffer2(458);	
			LineBuffer2(460) <= LineBuffer2(459);
			LineBuffer2(461) <= LineBuffer2(460);
			LineBuffer2(462) <= LineBuffer2(461);
			LineBuffer2(463) <= LineBuffer2(462);
			LineBuffer2(464) <= LineBuffer2(463);
			LineBuffer2(465) <= LineBuffer2(464);
			LineBuffer2(466) <= LineBuffer2(465);
			LineBuffer2(467) <= LineBuffer2(466);
			LineBuffer2(468) <= LineBuffer2(467);
			LineBuffer2(469) <= LineBuffer2(468);	
			LineBuffer2(470) <= LineBuffer2(469);
			LineBuffer2(471) <= LineBuffer2(470);
			LineBuffer2(472) <= LineBuffer2(471);
			LineBuffer2(473) <= LineBuffer2(472);
			LineBuffer2(474) <= LineBuffer2(473);
			LineBuffer2(475) <= LineBuffer2(474);
			LineBuffer2(476) <= LineBuffer2(475);
			LineBuffer2(477) <= LineBuffer2(476);
			LineBuffer2(478) <= LineBuffer2(477);
			LineBuffer2(479) <= LineBuffer2(478);	
			LineBuffer2(480) <= LineBuffer2(479);
			LineBuffer2(481) <= LineBuffer2(480);
			LineBuffer2(482) <= LineBuffer2(481);
			LineBuffer2(483) <= LineBuffer2(482);
			LineBuffer2(484) <= LineBuffer2(483);
			LineBuffer2(485) <= LineBuffer2(484);
			LineBuffer2(486) <= LineBuffer2(485);
			LineBuffer2(487) <= LineBuffer2(486);
			LineBuffer2(488) <= LineBuffer2(487);
			LineBuffer2(489) <= LineBuffer2(488);	
			LineBuffer2(490) <= LineBuffer2(489);
			LineBuffer2(491) <= LineBuffer2(490);
			LineBuffer2(492) <= LineBuffer2(491);
			LineBuffer2(493) <= LineBuffer2(492);
			LineBuffer2(494) <= LineBuffer2(493);
			LineBuffer2(495) <= LineBuffer2(494);
			LineBuffer2(496) <= LineBuffer2(495);
			LineBuffer2(497) <= LineBuffer2(496);
			LineBuffer2(498) <= LineBuffer2(497);
			LineBuffer2(499) <= LineBuffer2(498);	
			LineBuffer2(500) <= LineBuffer2(499);	
			LineBuffer2(501) <= LineBuffer2(500);
			LineBuffer2(502) <= LineBuffer2(501);
			LineBuffer2(503) <= LineBuffer2(502);
			LineBuffer2(504) <= LineBuffer2(503);
			LineBuffer2(505) <= LineBuffer2(504);
			LineBuffer2(506) <= LineBuffer2(505);
			LineBuffer2(507) <= LineBuffer2(506);
			LineBuffer2(508) <= LineBuffer2(507);
			LineBuffer2(509) <= LineBuffer2(508);	
			LineBuffer2(510) <= LineBuffer2(509);
			LineBuffer2(511) <= LineBuffer2(510);
			LineBuffer2(512) <= LineBuffer2(511);
			LineBuffer2(513) <= LineBuffer2(512);
			LineBuffer2(514) <= LineBuffer2(513);
			LineBuffer2(515) <= LineBuffer2(514);
			LineBuffer2(516) <= LineBuffer2(515);
			LineBuffer2(517) <= LineBuffer2(516);
			LineBuffer2(518) <= LineBuffer2(517);
			LineBuffer2(519) <= LineBuffer2(518);	
			LineBuffer2(520) <= LineBuffer2(519);
			LineBuffer2(521) <= LineBuffer2(520);
			LineBuffer2(522) <= LineBuffer2(521);
			LineBuffer2(523) <= LineBuffer2(522);
			LineBuffer2(524) <= LineBuffer2(523);
			LineBuffer2(525) <= LineBuffer2(524);
			LineBuffer2(526) <= LineBuffer2(525);
			LineBuffer2(527) <= LineBuffer2(526);
			LineBuffer2(528) <= LineBuffer2(527);
			LineBuffer2(529) <= LineBuffer2(528);	
			LineBuffer2(530) <= LineBuffer2(529);
			LineBuffer2(531) <= LineBuffer2(530);
			LineBuffer2(532) <= LineBuffer2(531);
			LineBuffer2(533) <= LineBuffer2(532);
			LineBuffer2(534) <= LineBuffer2(533);
			LineBuffer2(535) <= LineBuffer2(534);
			LineBuffer2(536) <= LineBuffer2(535);
			LineBuffer2(537) <= LineBuffer2(536);
			LineBuffer2(538) <= LineBuffer2(537);
			LineBuffer2(539) <= LineBuffer2(538);	
			LineBuffer2(540) <= LineBuffer2(539);
			LineBuffer2(541) <= LineBuffer2(540);
			LineBuffer2(542) <= LineBuffer2(541);
			LineBuffer2(543) <= LineBuffer2(542);
			LineBuffer2(544) <= LineBuffer2(543);
			LineBuffer2(545) <= LineBuffer2(544);
			LineBuffer2(546) <= LineBuffer2(545);
			LineBuffer2(547) <= LineBuffer2(546);
			LineBuffer2(548) <= LineBuffer2(547);
			LineBuffer2(549) <= LineBuffer2(548);	
			LineBuffer2(550) <= LineBuffer2(549);
			LineBuffer2(551) <= LineBuffer2(550);
			LineBuffer2(552) <= LineBuffer2(551);
			LineBuffer2(553) <= LineBuffer2(552);
			LineBuffer2(554) <= LineBuffer2(553);
			LineBuffer2(555) <= LineBuffer2(554);
			LineBuffer2(556) <= LineBuffer2(555);
			LineBuffer2(557) <= LineBuffer2(556);
			LineBuffer2(558) <= LineBuffer2(557);
			LineBuffer2(559) <= LineBuffer2(558);	
			LineBuffer2(560) <= LineBuffer2(559);
			LineBuffer2(561) <= LineBuffer2(560);
			LineBuffer2(562) <= LineBuffer2(561);
			LineBuffer2(563) <= LineBuffer2(562);
			LineBuffer2(564) <= LineBuffer2(563);
			LineBuffer2(565) <= LineBuffer2(564);
			LineBuffer2(566) <= LineBuffer2(565);
			LineBuffer2(567) <= LineBuffer2(566);
			LineBuffer2(568) <= LineBuffer2(567);
			LineBuffer2(569) <= LineBuffer2(568);	
			LineBuffer2(570) <= LineBuffer2(569);
			LineBuffer2(571) <= LineBuffer2(570);
			LineBuffer2(572) <= LineBuffer2(571);
			LineBuffer2(573) <= LineBuffer2(572);
			LineBuffer2(574) <= LineBuffer2(573);
			LineBuffer2(575) <= LineBuffer2(574);
			LineBuffer2(576) <= LineBuffer2(575);
			LineBuffer2(577) <= LineBuffer2(576);
			LineBuffer2(578) <= LineBuffer2(577);
			LineBuffer2(579) <= LineBuffer2(578);	
			LineBuffer2(580) <= LineBuffer2(579);
			LineBuffer2(581) <= LineBuffer2(580);
			LineBuffer2(582) <= LineBuffer2(581);
			LineBuffer2(583) <= LineBuffer2(582);
			LineBuffer2(584) <= LineBuffer2(583);
			LineBuffer2(585) <= LineBuffer2(584);
			LineBuffer2(586) <= LineBuffer2(585);
			LineBuffer2(587) <= LineBuffer2(586);
			LineBuffer2(588) <= LineBuffer2(587);
			LineBuffer2(589) <= LineBuffer2(588);	
			LineBuffer2(590) <= LineBuffer2(589);
			LineBuffer2(591) <= LineBuffer2(590);
			LineBuffer2(592) <= LineBuffer2(591);
			LineBuffer2(593) <= LineBuffer2(592);
			LineBuffer2(594) <= LineBuffer2(593);
			LineBuffer2(595) <= LineBuffer2(594);
			LineBuffer2(596) <= LineBuffer2(595);
			LineBuffer2(597) <= LineBuffer2(596);
			LineBuffer2(598) <= LineBuffer2(597);
			LineBuffer2(599) <= LineBuffer2(598);	
			LineBuffer2(600) <= LineBuffer2(599);	
			LineBuffer2(601) <= LineBuffer2(600);
			LineBuffer2(602) <= LineBuffer2(601);
			LineBuffer2(603) <= LineBuffer2(602);
			LineBuffer2(604) <= LineBuffer2(603);
			LineBuffer2(605) <= LineBuffer2(604);
			LineBuffer2(606) <= LineBuffer2(605);
			LineBuffer2(607) <= LineBuffer2(606);
			LineBuffer2(608) <= LineBuffer2(607);
			LineBuffer2(609) <= LineBuffer2(608);	
			LineBuffer2(610) <= LineBuffer2(609);
			LineBuffer2(611) <= LineBuffer2(610);
			LineBuffer2(612) <= LineBuffer2(611);
			LineBuffer2(613) <= LineBuffer2(612);
			LineBuffer2(614) <= LineBuffer2(613);
			LineBuffer2(615) <= LineBuffer2(614);
			LineBuffer2(616) <= LineBuffer2(615);
			LineBuffer2(617) <= LineBuffer2(616);
			LineBuffer2(618) <= LineBuffer2(617);
			LineBuffer2(619) <= LineBuffer2(618);	
			LineBuffer2(620) <= LineBuffer2(619);
			LineBuffer2(621) <= LineBuffer2(620);
			LineBuffer2(622) <= LineBuffer2(621);
			LineBuffer2(623) <= LineBuffer2(622);
			LineBuffer2(624) <= LineBuffer2(623);
			LineBuffer2(625) <= LineBuffer2(624);
			LineBuffer2(626) <= LineBuffer2(625);
			LineBuffer2(627) <= LineBuffer2(626);
			LineBuffer2(628) <= LineBuffer2(627);
			LineBuffer2(629) <= LineBuffer2(628);	
			LineBuffer2(630) <= LineBuffer2(629);
			LineBuffer2(631) <= LineBuffer2(630);
			LineBuffer2(632) <= LineBuffer2(631);
			LineBuffer2(633) <= LineBuffer2(632);
			LineBuffer2(634) <= LineBuffer2(633);
			LineBuffer2(635) <= LineBuffer2(634);
			LineBuffer2(636) <= LineBuffer2(635);
			LineBuffer2(637) <= LineBuffer2(636);
			LineBuffer2(638) <= LineBuffer2(637);
			LineBuffer2(639) <= LineBuffer2(638);
		    LineBuffer2(640) <= LineBuffer2(639);
            LineBuffer2(641) <= LineBuffer2(640);
            LineBuffer2(642) <= LineBuffer2(641);
            LineBuffer2(643) <= LineBuffer2(642);
            LineBuffer2(644) <= LineBuffer2(643);
            LineBuffer2(645) <= LineBuffer2(644);
            LineBuffer2(646) <= LineBuffer2(645);
            LineBuffer2(647) <= LineBuffer2(646);
            LineBuffer2(648) <= LineBuffer2(647);
            LineBuffer2(649) <= LineBuffer2(648);    
            LineBuffer2(650) <= LineBuffer2(649);
            LineBuffer2(651) <= LineBuffer2(650);
            LineBuffer2(652) <= LineBuffer2(651);
            LineBuffer2(653) <= LineBuffer2(652);
            LineBuffer2(654) <= LineBuffer2(653);
            LineBuffer2(655) <= LineBuffer2(654);
            LineBuffer2(656) <= LineBuffer2(655);
            LineBuffer2(657) <= LineBuffer2(656);
            LineBuffer2(658) <= LineBuffer2(657);
            LineBuffer2(659) <= LineBuffer2(658);    
            LineBuffer2(660) <= LineBuffer2(659);
            LineBuffer2(661) <= LineBuffer2(660);
            LineBuffer2(662) <= LineBuffer2(661);
            LineBuffer2(663) <= LineBuffer2(662);
            LineBuffer2(664) <= LineBuffer2(663);
            LineBuffer2(665) <= LineBuffer2(664);
            LineBuffer2(666) <= LineBuffer2(665);
            LineBuffer2(667) <= LineBuffer2(666);
            LineBuffer2(668) <= LineBuffer2(667);
            LineBuffer2(669) <= LineBuffer2(668);    
            LineBuffer2(670) <= LineBuffer2(669);
            LineBuffer2(671) <= LineBuffer2(670);
            LineBuffer2(672) <= LineBuffer2(671);
            LineBuffer2(673) <= LineBuffer2(672);
            LineBuffer2(674) <= LineBuffer2(673);
            LineBuffer2(675) <= LineBuffer2(674);
            LineBuffer2(676) <= LineBuffer2(675);
            LineBuffer2(677) <= LineBuffer2(676);
            LineBuffer2(678) <= LineBuffer2(677);
            LineBuffer2(679) <= LineBuffer2(678);    
            LineBuffer2(680) <= LineBuffer2(679);
            LineBuffer2(681) <= LineBuffer2(680);
            LineBuffer2(682) <= LineBuffer2(681);
            LineBuffer2(683) <= LineBuffer2(682);
            LineBuffer2(684) <= LineBuffer2(683);
            LineBuffer2(685) <= LineBuffer2(684);
            LineBuffer2(686) <= LineBuffer2(685);
            LineBuffer2(687) <= LineBuffer2(686);
            LineBuffer2(688) <= LineBuffer2(687);
            LineBuffer2(689) <= LineBuffer2(688);    
            LineBuffer2(690) <= LineBuffer2(689);
            LineBuffer2(691) <= LineBuffer2(690);
            LineBuffer2(692) <= LineBuffer2(691);
            LineBuffer2(693) <= LineBuffer2(692);
            LineBuffer2(694) <= LineBuffer2(693);
            LineBuffer2(695) <= LineBuffer2(694);
            LineBuffer2(696) <= LineBuffer2(695);
            LineBuffer2(697) <= LineBuffer2(696);
            LineBuffer2(698) <= LineBuffer2(697);
            LineBuffer2(699) <= LineBuffer2(698);    
            LineBuffer2(700) <= LineBuffer2(699);
            LineBuffer2(701) <= LineBuffer2(700);
            LineBuffer2(702) <= LineBuffer2(701);
            LineBuffer2(703) <= LineBuffer2(702);
            LineBuffer2(704) <= LineBuffer2(703);
            LineBuffer2(705) <= LineBuffer2(704);
            LineBuffer2(706) <= LineBuffer2(705);
            LineBuffer2(707) <= LineBuffer2(706);
            LineBuffer2(708) <= LineBuffer2(707);
            LineBuffer2(709) <= LineBuffer2(708);    
            LineBuffer2(710) <= LineBuffer2(709);
            LineBuffer2(711) <= LineBuffer2(710);
            LineBuffer2(712) <= LineBuffer2(711);
            LineBuffer2(713) <= LineBuffer2(712);
            LineBuffer2(714) <= LineBuffer2(713);
            LineBuffer2(715) <= LineBuffer2(714);
            LineBuffer2(716) <= LineBuffer2(715);
            LineBuffer2(717) <= LineBuffer2(716);
            LineBuffer2(718) <= LineBuffer2(717);
            LineBuffer2(719) <= LineBuffer2(718);    
            LineBuffer2(720) <= LineBuffer2(719);
            LineBuffer2(721) <= LineBuffer2(720);
            LineBuffer2(722) <= LineBuffer2(721);
            LineBuffer2(723) <= LineBuffer2(722);
            LineBuffer2(724) <= LineBuffer2(723);
            LineBuffer2(725) <= LineBuffer2(724);
            LineBuffer2(726) <= LineBuffer2(725);
            LineBuffer2(727) <= LineBuffer2(726);
            LineBuffer2(728) <= LineBuffer2(727);
            LineBuffer2(729) <= LineBuffer2(728);    
            LineBuffer2(730) <= LineBuffer2(729);
            LineBuffer2(731) <= LineBuffer2(730);
            LineBuffer2(732) <= LineBuffer2(731);
            LineBuffer2(733) <= LineBuffer2(732);
            LineBuffer2(734) <= LineBuffer2(733);
            LineBuffer2(735) <= LineBuffer2(734);
            LineBuffer2(736) <= LineBuffer2(735);
            LineBuffer2(737) <= LineBuffer2(736);
            LineBuffer2(738) <= LineBuffer2(737);
            LineBuffer2(739) <= LineBuffer2(738);    
            LineBuffer2(740) <= LineBuffer2(739);
            LineBuffer2(741) <= LineBuffer2(740);
            LineBuffer2(742) <= LineBuffer2(741);
            LineBuffer2(743) <= LineBuffer2(742);
            LineBuffer2(744) <= LineBuffer2(743);
            LineBuffer2(745) <= LineBuffer2(744);
            LineBuffer2(746) <= LineBuffer2(745);
            LineBuffer2(747) <= LineBuffer2(746);
            LineBuffer2(748) <= LineBuffer2(747);
            LineBuffer2(749) <= LineBuffer2(748);    
            LineBuffer2(750) <= LineBuffer2(749);
            LineBuffer2(751) <= LineBuffer2(750);
            LineBuffer2(752) <= LineBuffer2(751);
            LineBuffer2(753) <= LineBuffer2(752);
            LineBuffer2(754) <= LineBuffer2(753);
            LineBuffer2(755) <= LineBuffer2(754);
            LineBuffer2(756) <= LineBuffer2(755);
            LineBuffer2(757) <= LineBuffer2(756);
            LineBuffer2(758) <= LineBuffer2(757);
            LineBuffer2(759) <= LineBuffer2(758);    
            LineBuffer2(760) <= LineBuffer2(759);
            LineBuffer2(761) <= LineBuffer2(760);
            LineBuffer2(762) <= LineBuffer2(761);
            LineBuffer2(763) <= LineBuffer2(762);
            LineBuffer2(764) <= LineBuffer2(763);
            LineBuffer2(765) <= LineBuffer2(764);
            LineBuffer2(766) <= LineBuffer2(765);
            LineBuffer2(767) <= LineBuffer2(766);
            LineBuffer2(768) <= LineBuffer2(767);
            LineBuffer2(769) <= LineBuffer2(768);    
            LineBuffer2(770) <= LineBuffer2(769);
            LineBuffer2(771) <= LineBuffer2(770);
            LineBuffer2(772) <= LineBuffer2(771);
            LineBuffer2(773) <= LineBuffer2(772);
            LineBuffer2(774) <= LineBuffer2(773);
            LineBuffer2(775) <= LineBuffer2(774);
            LineBuffer2(776) <= LineBuffer2(775);
            LineBuffer2(777) <= LineBuffer2(776);
            LineBuffer2(778) <= LineBuffer2(777);
            LineBuffer2(779) <= LineBuffer2(778);    
            LineBuffer2(780) <= LineBuffer2(779);
            LineBuffer2(781) <= LineBuffer2(780);
            LineBuffer2(782) <= LineBuffer2(781);
            LineBuffer2(783) <= LineBuffer2(782);
            LineBuffer2(784) <= LineBuffer2(783);
            LineBuffer2(785) <= LineBuffer2(784);
            LineBuffer2(786) <= LineBuffer2(785);
            LineBuffer2(787) <= LineBuffer2(786);
            LineBuffer2(788) <= LineBuffer2(787);
            LineBuffer2(789) <= LineBuffer2(788);    
            LineBuffer2(790) <= LineBuffer2(789);
            LineBuffer2(791) <= LineBuffer2(790);
            LineBuffer2(792) <= LineBuffer2(791);
            LineBuffer2(793) <= LineBuffer2(792);
            LineBuffer2(794) <= LineBuffer2(793);
            LineBuffer2(795) <= LineBuffer2(794);
            LineBuffer2(796) <= LineBuffer2(795);
            LineBuffer2(797) <= LineBuffer2(796);
            LineBuffer2(798) <= LineBuffer2(797);
            LineBuffer2(799) <= LineBuffer2(798);    
            LineBuffer2(800) <= LineBuffer2(799);
            LineBuffer2(801) <= LineBuffer2(800);
            LineBuffer2(802) <= LineBuffer2(801);
            LineBuffer2(803) <= LineBuffer2(802);
            LineBuffer2(804) <= LineBuffer2(803);
            LineBuffer2(805) <= LineBuffer2(804);
            LineBuffer2(806) <= LineBuffer2(805);
            LineBuffer2(807) <= LineBuffer2(806);
            LineBuffer2(808) <= LineBuffer2(807);
            LineBuffer2(809) <= LineBuffer2(808);    
            LineBuffer2(810) <= LineBuffer2(809);
            LineBuffer2(811) <= LineBuffer2(810);
            LineBuffer2(812) <= LineBuffer2(811);
            LineBuffer2(813) <= LineBuffer2(812);
            LineBuffer2(814) <= LineBuffer2(813);
            LineBuffer2(815) <= LineBuffer2(814);
            LineBuffer2(816) <= LineBuffer2(815);
            LineBuffer2(817) <= LineBuffer2(816);
            LineBuffer2(818) <= LineBuffer2(817);
            LineBuffer2(819) <= LineBuffer2(818);    
            LineBuffer2(820) <= LineBuffer2(819);
            LineBuffer2(821) <= LineBuffer2(820);
            LineBuffer2(822) <= LineBuffer2(821);
            LineBuffer2(823) <= LineBuffer2(822);
            LineBuffer2(824) <= LineBuffer2(823);
            LineBuffer2(825) <= LineBuffer2(824);
            LineBuffer2(826) <= LineBuffer2(825);
            LineBuffer2(827) <= LineBuffer2(826);
            LineBuffer2(828) <= LineBuffer2(827);
            LineBuffer2(829) <= LineBuffer2(828);    
            LineBuffer2(830) <= LineBuffer2(829);
            LineBuffer2(831) <= LineBuffer2(830);
            LineBuffer2(832) <= LineBuffer2(831);
            LineBuffer2(833) <= LineBuffer2(832);
            LineBuffer2(834) <= LineBuffer2(833);
            LineBuffer2(835) <= LineBuffer2(834);
            LineBuffer2(836) <= LineBuffer2(835);
            LineBuffer2(837) <= LineBuffer2(836);
            LineBuffer2(838) <= LineBuffer2(837);
            LineBuffer2(839) <= LineBuffer2(838);
            LineBuffer2(840) <= LineBuffer2(839);
            LineBuffer2(841) <= LineBuffer2(840);
            LineBuffer2(842) <= LineBuffer2(841);
            LineBuffer2(843) <= LineBuffer2(842);
            LineBuffer2(844) <= LineBuffer2(843);
            LineBuffer2(845) <= LineBuffer2(844);
            LineBuffer2(846) <= LineBuffer2(845);
            LineBuffer2(847) <= LineBuffer2(846);
            LineBuffer2(848) <= LineBuffer2(847);
            LineBuffer2(849) <= LineBuffer2(848);    
            LineBuffer2(850) <= LineBuffer2(849);
            LineBuffer2(851) <= LineBuffer2(850);
            LineBuffer2(852) <= LineBuffer2(851);
            LineBuffer2(853) <= LineBuffer2(852);
            LineBuffer2(854) <= LineBuffer2(853);
            LineBuffer2(855) <= LineBuffer2(854);
            LineBuffer2(856) <= LineBuffer2(855);
            LineBuffer2(857) <= LineBuffer2(856);
            LineBuffer2(858) <= LineBuffer2(857);
            LineBuffer2(859) <= LineBuffer2(858);    
            LineBuffer2(860) <= LineBuffer2(859);
            LineBuffer2(861) <= LineBuffer2(860);
            LineBuffer2(862) <= LineBuffer2(861);
            LineBuffer2(863) <= LineBuffer2(862);
            LineBuffer2(864) <= LineBuffer2(863);
            LineBuffer2(865) <= LineBuffer2(864);
            LineBuffer2(866) <= LineBuffer2(865);
            LineBuffer2(867) <= LineBuffer2(866);
            LineBuffer2(868) <= LineBuffer2(867);
            LineBuffer2(869) <= LineBuffer2(868);    
            LineBuffer2(870) <= LineBuffer2(869);
            LineBuffer2(871) <= LineBuffer2(870);
            LineBuffer2(872) <= LineBuffer2(871);
            LineBuffer2(873) <= LineBuffer2(872);
            LineBuffer2(874) <= LineBuffer2(873);
            LineBuffer2(875) <= LineBuffer2(874);
            LineBuffer2(876) <= LineBuffer2(875);
            LineBuffer2(877) <= LineBuffer2(876);
            LineBuffer2(878) <= LineBuffer2(877);
            LineBuffer2(879) <= LineBuffer2(878);    
            LineBuffer2(880) <= LineBuffer2(879);
            LineBuffer2(881) <= LineBuffer2(880);
            LineBuffer2(882) <= LineBuffer2(881);
            LineBuffer2(883) <= LineBuffer2(882);
            LineBuffer2(884) <= LineBuffer2(883);
            LineBuffer2(885) <= LineBuffer2(884);
            LineBuffer2(886) <= LineBuffer2(885);
            LineBuffer2(887) <= LineBuffer2(886);
            LineBuffer2(888) <= LineBuffer2(887);
            LineBuffer2(889) <= LineBuffer2(888);    
            LineBuffer2(890) <= LineBuffer2(889);
            LineBuffer2(891) <= LineBuffer2(890);
            LineBuffer2(892) <= LineBuffer2(891);
            LineBuffer2(893) <= LineBuffer2(892);
            LineBuffer2(894) <= LineBuffer2(893);
            LineBuffer2(895) <= LineBuffer2(894);
            LineBuffer2(896) <= LineBuffer2(895);
            LineBuffer2(897) <= LineBuffer2(896);
            LineBuffer2(898) <= LineBuffer2(897);
            LineBuffer2(899) <= LineBuffer2(898);    
            LineBuffer2(900) <= LineBuffer2(899);
            LineBuffer2(901) <= LineBuffer2(900);
            LineBuffer2(902) <= LineBuffer2(901);
            LineBuffer2(903) <= LineBuffer2(902);
            LineBuffer2(904) <= LineBuffer2(903);
            LineBuffer2(905) <= LineBuffer2(904);
            LineBuffer2(906) <= LineBuffer2(905);
            LineBuffer2(907) <= LineBuffer2(906);
            LineBuffer2(908) <= LineBuffer2(907);
            LineBuffer2(909) <= LineBuffer2(908);    
            LineBuffer2(910) <= LineBuffer2(909);
            LineBuffer2(911) <= LineBuffer2(910);
            LineBuffer2(912) <= LineBuffer2(911);
            LineBuffer2(913) <= LineBuffer2(912);
            LineBuffer2(914) <= LineBuffer2(913);
            LineBuffer2(915) <= LineBuffer2(914);
            LineBuffer2(916) <= LineBuffer2(915);
            LineBuffer2(917) <= LineBuffer2(916);
            LineBuffer2(918) <= LineBuffer2(917);
            LineBuffer2(919) <= LineBuffer2(918);    
            LineBuffer2(920) <= LineBuffer2(919);
            LineBuffer2(921) <= LineBuffer2(920);
            LineBuffer2(922) <= LineBuffer2(921);
            LineBuffer2(923) <= LineBuffer2(922);
            LineBuffer2(924) <= LineBuffer2(923);
            LineBuffer2(925) <= LineBuffer2(924);
            LineBuffer2(926) <= LineBuffer2(925);
            LineBuffer2(927) <= LineBuffer2(926);
            LineBuffer2(928) <= LineBuffer2(927);
            LineBuffer2(929) <= LineBuffer2(928);    
            LineBuffer2(930) <= LineBuffer2(929);
            LineBuffer2(931) <= LineBuffer2(930);
            LineBuffer2(932) <= LineBuffer2(931);
            LineBuffer2(933) <= LineBuffer2(932);
            LineBuffer2(934) <= LineBuffer2(933);
            LineBuffer2(935) <= LineBuffer2(934);
            LineBuffer2(936) <= LineBuffer2(935);
            LineBuffer2(937) <= LineBuffer2(936);
            LineBuffer2(938) <= LineBuffer2(937);
            LineBuffer2(939) <= LineBuffer2(938);
            LineBuffer2(940) <= LineBuffer2(939);
            LineBuffer2(941) <= LineBuffer2(940);
            LineBuffer2(942) <= LineBuffer2(941);
            LineBuffer2(943) <= LineBuffer2(942);
            LineBuffer2(944) <= LineBuffer2(943);
            LineBuffer2(945) <= LineBuffer2(944);
            LineBuffer2(946) <= LineBuffer2(945);
            LineBuffer2(947) <= LineBuffer2(946);
            LineBuffer2(948) <= LineBuffer2(947);
            LineBuffer2(949) <= LineBuffer2(948);    
            LineBuffer2(950) <= LineBuffer2(949);
            LineBuffer2(951) <= LineBuffer2(950);
            LineBuffer2(952) <= LineBuffer2(951);
            LineBuffer2(953) <= LineBuffer2(952);
            LineBuffer2(954) <= LineBuffer2(953);
            LineBuffer2(955) <= LineBuffer2(954);
            LineBuffer2(956) <= LineBuffer2(955);
            LineBuffer2(957) <= LineBuffer2(956);
            LineBuffer2(958) <= LineBuffer2(957);
            LineBuffer2(959) <= LineBuffer2(958);    
            LineBuffer2(960) <= LineBuffer2(959);
            LineBuffer2(961) <= LineBuffer2(960);
            LineBuffer2(962) <= LineBuffer2(961);
            LineBuffer2(963) <= LineBuffer2(962);
            LineBuffer2(964) <= LineBuffer2(963);
            LineBuffer2(965) <= LineBuffer2(964);
            LineBuffer2(966) <= LineBuffer2(965);
            LineBuffer2(967) <= LineBuffer2(966);
            LineBuffer2(968) <= LineBuffer2(967);
            LineBuffer2(969) <= LineBuffer2(968);    
            LineBuffer2(970) <= LineBuffer2(969);
            LineBuffer2(971) <= LineBuffer2(970);
            LineBuffer2(972) <= LineBuffer2(971);
            LineBuffer2(973) <= LineBuffer2(972);
            LineBuffer2(974) <= LineBuffer2(973);
            LineBuffer2(975) <= LineBuffer2(974);
            LineBuffer2(976) <= LineBuffer2(975);
            LineBuffer2(977) <= LineBuffer2(976);
            LineBuffer2(978) <= LineBuffer2(977);
            LineBuffer2(979) <= LineBuffer2(978);    
            LineBuffer2(980) <= LineBuffer2(979);
            LineBuffer2(981) <= LineBuffer2(980);
            LineBuffer2(982) <= LineBuffer2(981);
            LineBuffer2(983) <= LineBuffer2(982);
            LineBuffer2(984) <= LineBuffer2(983);
            LineBuffer2(985) <= LineBuffer2(984);
            LineBuffer2(986) <= LineBuffer2(985);
            LineBuffer2(987) <= LineBuffer2(986);
            LineBuffer2(988) <= LineBuffer2(987);
            LineBuffer2(989) <= LineBuffer2(988);    
            LineBuffer2(990) <= LineBuffer2(989);
            LineBuffer2(991) <= LineBuffer2(990);
            LineBuffer2(992) <= LineBuffer2(991);
            LineBuffer2(993) <= LineBuffer2(992);
            LineBuffer2(994) <= LineBuffer2(993);
            LineBuffer2(995) <= LineBuffer2(994);
            LineBuffer2(996) <= LineBuffer2(995);
            LineBuffer2(997) <= LineBuffer2(996);
            LineBuffer2(998) <= LineBuffer2(997);
            LineBuffer2(999) <= LineBuffer2(998);    
            LineBuffer2(1000) <= LineBuffer2(999);
            LineBuffer2(1001) <= LineBuffer2(1000);
            LineBuffer2(1002) <= LineBuffer2(1001);
            LineBuffer2(1003) <= LineBuffer2(1002);
            LineBuffer2(1004) <= LineBuffer2(1003);
            LineBuffer2(1005) <= LineBuffer2(1004);
            LineBuffer2(1006) <= LineBuffer2(1005);
            LineBuffer2(1007) <= LineBuffer2(1006);
            LineBuffer2(1008) <= LineBuffer2(1007);
            LineBuffer2(1009) <= LineBuffer2(1008);    
            LineBuffer2(1010) <= LineBuffer2(1009);
            LineBuffer2(1011) <= LineBuffer2(1010);
            LineBuffer2(1012) <= LineBuffer2(1011);
            LineBuffer2(1013) <= LineBuffer2(1012);
            LineBuffer2(1014) <= LineBuffer2(1013);
            LineBuffer2(1015) <= LineBuffer2(1014);
            LineBuffer2(1016) <= LineBuffer2(1015);
            LineBuffer2(1017) <= LineBuffer2(1016);
            LineBuffer2(1018) <= LineBuffer2(1017);
            LineBuffer2(1019) <= LineBuffer2(1018);    
            LineBuffer2(1020) <= LineBuffer2(1019);
            LineBuffer2(1021) <= LineBuffer2(1020);
            LineBuffer2(1022) <= LineBuffer2(1021);
            LineBuffer2(1023) <= LineBuffer2(1022);
            LineBuffer2(1024) <= LineBuffer2(1023);
            LineBuffer2(1025) <= LineBuffer2(1024);
            LineBuffer2(1026) <= LineBuffer2(1025);
            LineBuffer2(1027) <= LineBuffer2(1026);
            LineBuffer2(1028) <= LineBuffer2(1027);
            LineBuffer2(1029) <= LineBuffer2(1028);    
            LineBuffer2(1030) <= LineBuffer2(1029);
            LineBuffer2(1031) <= LineBuffer2(1030);
            LineBuffer2(1032) <= LineBuffer2(1031);
            LineBuffer2(1033) <= LineBuffer2(1032);
            LineBuffer2(1034) <= LineBuffer2(1033);
            LineBuffer2(1035) <= LineBuffer2(1034);
            LineBuffer2(1036) <= LineBuffer2(1035);
            LineBuffer2(1037) <= LineBuffer2(1036);
            LineBuffer2(1038) <= LineBuffer2(1037);
            LineBuffer2(1039) <= LineBuffer2(1038);
            LineBuffer2(1040) <= LineBuffer2(1039);
            LineBuffer2(1041) <= LineBuffer2(1040);
            LineBuffer2(1042) <= LineBuffer2(1041);
            LineBuffer2(1043) <= LineBuffer2(1042);
            LineBuffer2(1044) <= LineBuffer2(1043);
            LineBuffer2(1045) <= LineBuffer2(1044);
            LineBuffer2(1046) <= LineBuffer2(1045);
            LineBuffer2(1047) <= LineBuffer2(1046);
            LineBuffer2(1048) <= LineBuffer2(1047);
            LineBuffer2(1049) <= LineBuffer2(1048);    
            LineBuffer2(1050) <= LineBuffer2(1049);
            LineBuffer2(1051) <= LineBuffer2(1050);
            LineBuffer2(1052) <= LineBuffer2(1051);
            LineBuffer2(1053) <= LineBuffer2(1052);
            LineBuffer2(1054) <= LineBuffer2(1053);
            LineBuffer2(1055) <= LineBuffer2(1054);
            LineBuffer2(1056) <= LineBuffer2(1055);
            LineBuffer2(1057) <= LineBuffer2(1056);
            LineBuffer2(1058) <= LineBuffer2(1057);
            LineBuffer2(1059) <= LineBuffer2(1058);    
            LineBuffer2(1060) <= LineBuffer2(1059);
            LineBuffer2(1061) <= LineBuffer2(1060);
            LineBuffer2(1062) <= LineBuffer2(1061);
            LineBuffer2(1063) <= LineBuffer2(1062);
            LineBuffer2(1064) <= LineBuffer2(1063);
            LineBuffer2(1065) <= LineBuffer2(1064);
            LineBuffer2(1066) <= LineBuffer2(1065);
            LineBuffer2(1067) <= LineBuffer2(1066);
            LineBuffer2(1068) <= LineBuffer2(1067);
            LineBuffer2(1069) <= LineBuffer2(1068);    
            LineBuffer2(1070) <= LineBuffer2(1069);
            LineBuffer2(1071) <= LineBuffer2(1070);
            LineBuffer2(1072) <= LineBuffer2(1071);
            LineBuffer2(1073) <= LineBuffer2(1072);
            LineBuffer2(1074) <= LineBuffer2(1073);
            LineBuffer2(1075) <= LineBuffer2(1074);
            LineBuffer2(1076) <= LineBuffer2(1075);
            LineBuffer2(1077) <= LineBuffer2(1076);
            LineBuffer2(1078) <= LineBuffer2(1077);
            LineBuffer2(1079) <= LineBuffer2(1078);    
            LineBuffer2(1080) <= LineBuffer2(1079);
            LineBuffer2(1081) <= LineBuffer2(1080);
            LineBuffer2(1082) <= LineBuffer2(1081);
            LineBuffer2(1083) <= LineBuffer2(1082);
            LineBuffer2(1084) <= LineBuffer2(1083);
            LineBuffer2(1085) <= LineBuffer2(1084);
            LineBuffer2(1086) <= LineBuffer2(1085);
            LineBuffer2(1087) <= LineBuffer2(1086);
            LineBuffer2(1088) <= LineBuffer2(1087);
            LineBuffer2(1089) <= LineBuffer2(1088);    
            LineBuffer2(1090) <= LineBuffer2(1089);
            LineBuffer2(1091) <= LineBuffer2(1090);
            LineBuffer2(1092) <= LineBuffer2(1091);
            LineBuffer2(1093) <= LineBuffer2(1092);
            LineBuffer2(1094) <= LineBuffer2(1093);
            LineBuffer2(1095) <= LineBuffer2(1094);
            LineBuffer2(1096) <= LineBuffer2(1095);
            LineBuffer2(1097) <= LineBuffer2(1096);
            LineBuffer2(1098) <= LineBuffer2(1097);
            LineBuffer2(1099) <= LineBuffer2(1098);    
            LineBuffer2(1100) <= LineBuffer2(1099);
            LineBuffer2(1101) <= LineBuffer2(1100);
            LineBuffer2(1102) <= LineBuffer2(1101);
            LineBuffer2(1103) <= LineBuffer2(1102);
            LineBuffer2(1104) <= LineBuffer2(1103);
            LineBuffer2(1105) <= LineBuffer2(1104);
            LineBuffer2(1106) <= LineBuffer2(1105);
            LineBuffer2(1107) <= LineBuffer2(1106);
            LineBuffer2(1108) <= LineBuffer2(1107);
            LineBuffer2(1109) <= LineBuffer2(1108);    
            LineBuffer2(1110) <= LineBuffer2(1109);
            LineBuffer2(1111) <= LineBuffer2(1110);
            LineBuffer2(1112) <= LineBuffer2(1111);
            LineBuffer2(1113) <= LineBuffer2(1112);
            LineBuffer2(1114) <= LineBuffer2(1113);
            LineBuffer2(1115) <= LineBuffer2(1114);
            LineBuffer2(1116) <= LineBuffer2(1115);
            LineBuffer2(1117) <= LineBuffer2(1116);
            LineBuffer2(1118) <= LineBuffer2(1117);
            LineBuffer2(1119) <= LineBuffer2(1118);    
            LineBuffer2(1120) <= LineBuffer2(1119);
            LineBuffer2(1121) <= LineBuffer2(1120);
            LineBuffer2(1122) <= LineBuffer2(1121);
            LineBuffer2(1123) <= LineBuffer2(1122);
            LineBuffer2(1124) <= LineBuffer2(1123);
            LineBuffer2(1125) <= LineBuffer2(1124);
            LineBuffer2(1126) <= LineBuffer2(1125);
            LineBuffer2(1127) <= LineBuffer2(1126);
            LineBuffer2(1128) <= LineBuffer2(1127);
            LineBuffer2(1129) <= LineBuffer2(1128);    
            LineBuffer2(1130) <= LineBuffer2(1129);
            LineBuffer2(1131) <= LineBuffer2(1130);
            LineBuffer2(1132) <= LineBuffer2(1131);
            LineBuffer2(1133) <= LineBuffer2(1132);
            LineBuffer2(1134) <= LineBuffer2(1133);
            LineBuffer2(1135) <= LineBuffer2(1134);
            LineBuffer2(1136) <= LineBuffer2(1135);
            LineBuffer2(1137) <= LineBuffer2(1136);
            LineBuffer2(1138) <= LineBuffer2(1137);
            LineBuffer2(1139) <= LineBuffer2(1138);
            LineBuffer2(1140) <= LineBuffer2(1139);
            LineBuffer2(1141) <= LineBuffer2(1140);
            LineBuffer2(1142) <= LineBuffer2(1141);
            LineBuffer2(1143) <= LineBuffer2(1142);
            LineBuffer2(1144) <= LineBuffer2(1143);
            LineBuffer2(1145) <= LineBuffer2(1144);
            LineBuffer2(1146) <= LineBuffer2(1145);
            LineBuffer2(1147) <= LineBuffer2(1146);
            LineBuffer2(1148) <= LineBuffer2(1147);
            LineBuffer2(1149) <= LineBuffer2(1148);    
            LineBuffer2(1150) <= LineBuffer2(1149);
            LineBuffer2(1151) <= LineBuffer2(1150);
            LineBuffer2(1152) <= LineBuffer2(1151);
            LineBuffer2(1153) <= LineBuffer2(1152);
            LineBuffer2(1154) <= LineBuffer2(1153);
            LineBuffer2(1155) <= LineBuffer2(1154);
            LineBuffer2(1156) <= LineBuffer2(1155);
            LineBuffer2(1157) <= LineBuffer2(1156);
            LineBuffer2(1158) <= LineBuffer2(1157);
            LineBuffer2(1159) <= LineBuffer2(1158);    
            LineBuffer2(1160) <= LineBuffer2(1159);
            LineBuffer2(1161) <= LineBuffer2(1160);
            LineBuffer2(1162) <= LineBuffer2(1161);
            LineBuffer2(1163) <= LineBuffer2(1162);
            LineBuffer2(1164) <= LineBuffer2(1163);
            LineBuffer2(1165) <= LineBuffer2(1164);
            LineBuffer2(1166) <= LineBuffer2(1165);
            LineBuffer2(1167) <= LineBuffer2(1166);
            LineBuffer2(1168) <= LineBuffer2(1167);
            LineBuffer2(1169) <= LineBuffer2(1168);    
            LineBuffer2(1170) <= LineBuffer2(1169);
            LineBuffer2(1171) <= LineBuffer2(1170);
            LineBuffer2(1172) <= LineBuffer2(1171);
            LineBuffer2(1173) <= LineBuffer2(1172);
            LineBuffer2(1174) <= LineBuffer2(1173);
            LineBuffer2(1175) <= LineBuffer2(1174);
            LineBuffer2(1176) <= LineBuffer2(1175);
            LineBuffer2(1177) <= LineBuffer2(1176);
            LineBuffer2(1178) <= LineBuffer2(1177);
            LineBuffer2(1179) <= LineBuffer2(1178);    
            LineBuffer2(1180) <= LineBuffer2(1179);
            LineBuffer2(1181) <= LineBuffer2(1180);
            LineBuffer2(1182) <= LineBuffer2(1181);
            LineBuffer2(1183) <= LineBuffer2(1182);
            LineBuffer2(1184) <= LineBuffer2(1183);
            LineBuffer2(1185) <= LineBuffer2(1184);
            LineBuffer2(1186) <= LineBuffer2(1185);
            LineBuffer2(1187) <= LineBuffer2(1186);
            LineBuffer2(1188) <= LineBuffer2(1187);
            LineBuffer2(1189) <= LineBuffer2(1188);    
            LineBuffer2(1190) <= LineBuffer2(1189);
            LineBuffer2(1191) <= LineBuffer2(1190);
            LineBuffer2(1192) <= LineBuffer2(1191);
            LineBuffer2(1193) <= LineBuffer2(1192);
            LineBuffer2(1194) <= LineBuffer2(1193);
            LineBuffer2(1195) <= LineBuffer2(1194);
            LineBuffer2(1196) <= LineBuffer2(1195);
            LineBuffer2(1197) <= LineBuffer2(1196);
            LineBuffer2(1198) <= LineBuffer2(1197);
            LineBuffer2(1199) <= LineBuffer2(1198);    
            LineBuffer2(1200) <= LineBuffer2(1199);
            LineBuffer2(1201) <= LineBuffer2(1200);
            LineBuffer2(1202) <= LineBuffer2(1201);
            LineBuffer2(1203) <= LineBuffer2(1202);
            LineBuffer2(1204) <= LineBuffer2(1203);
            LineBuffer2(1205) <= LineBuffer2(1204);
            LineBuffer2(1206) <= LineBuffer2(1205);
            LineBuffer2(1207) <= LineBuffer2(1206);
            LineBuffer2(1208) <= LineBuffer2(1207);
            LineBuffer2(1209) <= LineBuffer2(1208);    
            LineBuffer2(1210) <= LineBuffer2(1209);
            LineBuffer2(1211) <= LineBuffer2(1210);
            LineBuffer2(1212) <= LineBuffer2(1211);
            LineBuffer2(1213) <= LineBuffer2(1212);
            LineBuffer2(1214) <= LineBuffer2(1213);
            LineBuffer2(1215) <= LineBuffer2(1214);
            LineBuffer2(1216) <= LineBuffer2(1215);
            LineBuffer2(1217) <= LineBuffer2(1216);
            LineBuffer2(1218) <= LineBuffer2(1217);
            LineBuffer2(1219) <= LineBuffer2(1218);    
            LineBuffer2(1220) <= LineBuffer2(1219);
            LineBuffer2(1221) <= LineBuffer2(1220);
            LineBuffer2(1222) <= LineBuffer2(1221);
            LineBuffer2(1223) <= LineBuffer2(1222);
            LineBuffer2(1224) <= LineBuffer2(1223);
            LineBuffer2(1225) <= LineBuffer2(1224);
            LineBuffer2(1226) <= LineBuffer2(1225);
            LineBuffer2(1227) <= LineBuffer2(1226);
            LineBuffer2(1228) <= LineBuffer2(1227);
            LineBuffer2(1229) <= LineBuffer2(1228);    
            LineBuffer2(1230) <= LineBuffer2(1229);
            LineBuffer2(1231) <= LineBuffer2(1230);
            LineBuffer2(1232) <= LineBuffer2(1231);
            LineBuffer2(1233) <= LineBuffer2(1232);
            LineBuffer2(1234) <= LineBuffer2(1233);
            LineBuffer2(1235) <= LineBuffer2(1234);
            LineBuffer2(1236) <= LineBuffer2(1235);
            LineBuffer2(1237) <= LineBuffer2(1236);
            LineBuffer2(1238) <= LineBuffer2(1237);
            LineBuffer2(1239) <= LineBuffer2(1238);
            LineBuffer2(1240) <= LineBuffer2(1239);
            LineBuffer2(1241) <= LineBuffer2(1240);
            LineBuffer2(1242) <= LineBuffer2(1241);
            LineBuffer2(1243) <= LineBuffer2(1242);
            LineBuffer2(1244) <= LineBuffer2(1243);
            LineBuffer2(1245) <= LineBuffer2(1244);
            LineBuffer2(1246) <= LineBuffer2(1245);
            LineBuffer2(1247) <= LineBuffer2(1246);
            LineBuffer2(1248) <= LineBuffer2(1247);
            LineBuffer2(1249) <= LineBuffer2(1248);    
            LineBuffer2(1250) <= LineBuffer2(1249);
            LineBuffer2(1251) <= LineBuffer2(1250);
            LineBuffer2(1252) <= LineBuffer2(1251);
            LineBuffer2(1253) <= LineBuffer2(1252);
            LineBuffer2(1254) <= LineBuffer2(1253);
            LineBuffer2(1255) <= LineBuffer2(1254);
            LineBuffer2(1256) <= LineBuffer2(1255);
            LineBuffer2(1257) <= LineBuffer2(1256);
            LineBuffer2(1258) <= LineBuffer2(1257);
            LineBuffer2(1259) <= LineBuffer2(1258);    
            LineBuffer2(1260) <= LineBuffer2(1259);
            LineBuffer2(1261) <= LineBuffer2(1260);
            LineBuffer2(1262) <= LineBuffer2(1261);
            LineBuffer2(1263) <= LineBuffer2(1262);
            LineBuffer2(1264) <= LineBuffer2(1263);
            LineBuffer2(1265) <= LineBuffer2(1264);
            LineBuffer2(1266) <= LineBuffer2(1265);
            LineBuffer2(1267) <= LineBuffer2(1266);
            LineBuffer2(1268) <= LineBuffer2(1267);
            LineBuffer2(1269) <= LineBuffer2(1268);    
            LineBuffer2(1270) <= LineBuffer2(1269);
            LineBuffer2(1271) <= LineBuffer2(1270);
            LineBuffer2(1272) <= LineBuffer2(1271);
            LineBuffer2(1273) <= LineBuffer2(1272);
            LineBuffer2(1274) <= LineBuffer2(1273);
            LineBuffer2(1275) <= LineBuffer2(1274);
            LineBuffer2(1276) <= LineBuffer2(1275);
            LineBuffer2(1277) <= LineBuffer2(1276);
            LineBuffer2(1278) <= LineBuffer2(1277);
            LineBuffer2(1279) <= LineBuffer2(1278);
--            LineBuffer2(1280) <= LineBuffer2(1279);
--            LineBuffer2(1281) <= LineBuffer2(1280);
--            LineBuffer2(1282) <= LineBuffer2(1281);
--            LineBuffer2(1283) <= LineBuffer2(1282);
--            LineBuffer2(1284) <= LineBuffer2(1283);
--            LineBuffer2(1285) <= LineBuffer2(1284);
--            LineBuffer2(1286) <= LineBuffer2(1285);
--            LineBuffer2(1287) <= LineBuffer2(1286);
--            LineBuffer2(1288) <= LineBuffer2(1287);
--            LineBuffer2(1289) <= LineBuffer2(1288);    
--            LineBuffer2(1290) <= LineBuffer2(1289);
--            LineBuffer2(1291) <= LineBuffer2(1290);
--            LineBuffer2(1292) <= LineBuffer2(1291);
--            LineBuffer2(1293) <= LineBuffer2(1292);
--            LineBuffer2(1294) <= LineBuffer2(1293);
--            LineBuffer2(1295) <= LineBuffer2(1294);
--            LineBuffer2(1296) <= LineBuffer2(1295);
--            LineBuffer2(1297) <= LineBuffer2(1296);
--            LineBuffer2(1298) <= LineBuffer2(1297);
--            LineBuffer2(1299) <= LineBuffer2(1298);    
--            LineBuffer2(1300) <= LineBuffer2(1299);
--            LineBuffer2(1301) <= LineBuffer2(1300);
--            LineBuffer2(1302) <= LineBuffer2(1301);
--            LineBuffer2(1303) <= LineBuffer2(1302);
--            LineBuffer2(1304) <= LineBuffer2(1303);
--            LineBuffer2(1305) <= LineBuffer2(1304);
--            LineBuffer2(1306) <= LineBuffer2(1305);
--            LineBuffer2(1307) <= LineBuffer2(1306);
--            LineBuffer2(1308) <= LineBuffer2(1307);
--            LineBuffer2(1309) <= LineBuffer2(1308);    
--            LineBuffer2(1310) <= LineBuffer2(1309);
--            LineBuffer2(1311) <= LineBuffer2(1310);
--            LineBuffer2(1312) <= LineBuffer2(1311);
--            LineBuffer2(1313) <= LineBuffer2(1312);
--            LineBuffer2(1314) <= LineBuffer2(1313);
--            LineBuffer2(1315) <= LineBuffer2(1314);
--            LineBuffer2(1316) <= LineBuffer2(1315);
--            LineBuffer2(1317) <= LineBuffer2(1316);
--            LineBuffer2(1318) <= LineBuffer2(1317);
--            LineBuffer2(1319) <= LineBuffer2(1318);    
--            LineBuffer2(1320) <= LineBuffer2(1319);
--            LineBuffer2(1321) <= LineBuffer2(1320);
--            LineBuffer2(1322) <= LineBuffer2(1321);
--            LineBuffer2(1323) <= LineBuffer2(1322);
--            LineBuffer2(1324) <= LineBuffer2(1323);
--            LineBuffer2(1325) <= LineBuffer2(1324);
--            LineBuffer2(1326) <= LineBuffer2(1325);
--            LineBuffer2(1327) <= LineBuffer2(1326);
--            LineBuffer2(1328) <= LineBuffer2(1327);
--            LineBuffer2(1329) <= LineBuffer2(1328);    
--            LineBuffer2(1330) <= LineBuffer2(1329);
--            LineBuffer2(1331) <= LineBuffer2(1330);
--            LineBuffer2(1332) <= LineBuffer2(1331);
--            LineBuffer2(1333) <= LineBuffer2(1332);
--            LineBuffer2(1334) <= LineBuffer2(1333);
--            LineBuffer2(1335) <= LineBuffer2(1334);
--            LineBuffer2(1336) <= LineBuffer2(1335);
--            LineBuffer2(1337) <= LineBuffer2(1336);
--            LineBuffer2(1338) <= LineBuffer2(1337);
--            LineBuffer2(1339) <= LineBuffer2(1338);    
--            LineBuffer2(1340) <= LineBuffer2(1339);
--            LineBuffer2(1341) <= LineBuffer2(1340);
--            LineBuffer2(1342) <= LineBuffer2(1341);
--            LineBuffer2(1343) <= LineBuffer2(1342);
--            LineBuffer2(1344) <= LineBuffer2(1343);
--            LineBuffer2(1345) <= LineBuffer2(1344);
--            LineBuffer2(1346) <= LineBuffer2(1345);
--            LineBuffer2(1347) <= LineBuffer2(1346);
--            LineBuffer2(1348) <= LineBuffer2(1347);
--            LineBuffer2(1349) <= LineBuffer2(1348);    
--            LineBuffer2(1350) <= LineBuffer2(1349);
--            LineBuffer2(1351) <= LineBuffer2(1350);
--            LineBuffer2(1352) <= LineBuffer2(1351);
--            LineBuffer2(1353) <= LineBuffer2(1352);
--            LineBuffer2(1354) <= LineBuffer2(1353);
--            LineBuffer2(1355) <= LineBuffer2(1354);
--            LineBuffer2(1356) <= LineBuffer2(1355);
--            LineBuffer2(1357) <= LineBuffer2(1356);
--            LineBuffer2(1358) <= LineBuffer2(1357);
--            LineBuffer2(1359) <= LineBuffer2(1358);    
--            LineBuffer2(1360) <= LineBuffer2(1359);
--            LineBuffer2(1361) <= LineBuffer2(1360);
--            LineBuffer2(1362) <= LineBuffer2(1361);
--            LineBuffer2(1363) <= LineBuffer2(1362);
--            LineBuffer2(1364) <= LineBuffer2(1363);
--            LineBuffer2(1365) <= LineBuffer2(1364);
--            LineBuffer2(1366) <= LineBuffer2(1365);
--            LineBuffer2(1367) <= LineBuffer2(1366);
--            LineBuffer2(1368) <= LineBuffer2(1367);
--            LineBuffer2(1369) <= LineBuffer2(1368);    
--            LineBuffer2(1370) <= LineBuffer2(1369);
--            LineBuffer2(1371) <= LineBuffer2(1370);
--            LineBuffer2(1372) <= LineBuffer2(1371);
--            LineBuffer2(1373) <= LineBuffer2(1372);
--            LineBuffer2(1374) <= LineBuffer2(1373);
--            LineBuffer2(1375) <= LineBuffer2(1374);
--            LineBuffer2(1376) <= LineBuffer2(1375);
--            LineBuffer2(1377) <= LineBuffer2(1376);
--            LineBuffer2(1378) <= LineBuffer2(1377);
--            LineBuffer2(1379) <= LineBuffer2(1378);    
--            LineBuffer2(1380) <= LineBuffer2(1379);
--            LineBuffer2(1381) <= LineBuffer2(1380);
--            LineBuffer2(1382) <= LineBuffer2(1381);
--            LineBuffer2(1383) <= LineBuffer2(1382);
--            LineBuffer2(1384) <= LineBuffer2(1383);
--            LineBuffer2(1385) <= LineBuffer2(1384);
--            LineBuffer2(1386) <= LineBuffer2(1385);
--            LineBuffer2(1387) <= LineBuffer2(1386);
--            LineBuffer2(1388) <= LineBuffer2(1387);
--            LineBuffer2(1389) <= LineBuffer2(1388);    
--            LineBuffer2(1390) <= LineBuffer2(1389);
--            LineBuffer2(1391) <= LineBuffer2(1390);
--            LineBuffer2(1392) <= LineBuffer2(1391);
--            LineBuffer2(1393) <= LineBuffer2(1392);
--            LineBuffer2(1394) <= LineBuffer2(1393);
--            LineBuffer2(1395) <= LineBuffer2(1394);
--            LineBuffer2(1396) <= LineBuffer2(1395);
--            LineBuffer2(1397) <= LineBuffer2(1396);
--            LineBuffer2(1398) <= LineBuffer2(1397);
--            LineBuffer2(1399) <= LineBuffer2(1398);    
--            LineBuffer2(1400) <= LineBuffer2(1399);
--            LineBuffer2(1401) <= LineBuffer2(1400);
--            LineBuffer2(1402) <= LineBuffer2(1401);
--            LineBuffer2(1403) <= LineBuffer2(1402);
--            LineBuffer2(1404) <= LineBuffer2(1403);
--            LineBuffer2(1405) <= LineBuffer2(1404);
--            LineBuffer2(1406) <= LineBuffer2(1405);
--            LineBuffer2(1407) <= LineBuffer2(1406);
--            LineBuffer2(1408) <= LineBuffer2(1407);
--            LineBuffer2(1409) <= LineBuffer2(1408);    
--            LineBuffer2(1410) <= LineBuffer2(1409);
--            LineBuffer2(1411) <= LineBuffer2(1410);
--            LineBuffer2(1412) <= LineBuffer2(1411);
--            LineBuffer2(1413) <= LineBuffer2(1412);
--            LineBuffer2(1414) <= LineBuffer2(1413);
--            LineBuffer2(1415) <= LineBuffer2(1414);
--            LineBuffer2(1416) <= LineBuffer2(1415);
--            LineBuffer2(1417) <= LineBuffer2(1416);
--            LineBuffer2(1418) <= LineBuffer2(1417);
--            LineBuffer2(1419) <= LineBuffer2(1418);    
--            LineBuffer2(1420) <= LineBuffer2(1419);
--            LineBuffer2(1421) <= LineBuffer2(1420);
--            LineBuffer2(1422) <= LineBuffer2(1421);
--            LineBuffer2(1423) <= LineBuffer2(1422);
--            LineBuffer2(1424) <= LineBuffer2(1423);
--            LineBuffer2(1425) <= LineBuffer2(1424);
--            LineBuffer2(1426) <= LineBuffer2(1425);
--            LineBuffer2(1427) <= LineBuffer2(1426);
--            LineBuffer2(1428) <= LineBuffer2(1427);
--            LineBuffer2(1429) <= LineBuffer2(1428);    
--            LineBuffer2(1430) <= LineBuffer2(1429);
--            LineBuffer2(1431) <= LineBuffer2(1430);
--            LineBuffer2(1432) <= LineBuffer2(1431);
--            LineBuffer2(1433) <= LineBuffer2(1432);
--            LineBuffer2(1434) <= LineBuffer2(1433);
--            LineBuffer2(1435) <= LineBuffer2(1434);
--            LineBuffer2(1436) <= LineBuffer2(1435);
--            LineBuffer2(1437) <= LineBuffer2(1436);
--            LineBuffer2(1438) <= LineBuffer2(1437);
--            LineBuffer2(1439) <= LineBuffer2(1438);    
--            LineBuffer2(1440) <= LineBuffer2(1439);
--            LineBuffer2(1441) <= LineBuffer2(1440);
--            LineBuffer2(1442) <= LineBuffer2(1441);
--            LineBuffer2(1443) <= LineBuffer2(1442);
--            LineBuffer2(1444) <= LineBuffer2(1443);
--            LineBuffer2(1445) <= LineBuffer2(1444);
--            LineBuffer2(1446) <= LineBuffer2(1445);
--            LineBuffer2(1447) <= LineBuffer2(1446);
--            LineBuffer2(1448) <= LineBuffer2(1447);
--            LineBuffer2(1449) <= LineBuffer2(1448);    
--            LineBuffer2(1450) <= LineBuffer2(1449);
--            LineBuffer2(1451) <= LineBuffer2(1450);
--            LineBuffer2(1452) <= LineBuffer2(1451);
--            LineBuffer2(1453) <= LineBuffer2(1452);
--            LineBuffer2(1454) <= LineBuffer2(1453);
--            LineBuffer2(1455) <= LineBuffer2(1454);
--            LineBuffer2(1456) <= LineBuffer2(1455);
--            LineBuffer2(1457) <= LineBuffer2(1456);
--            LineBuffer2(1458) <= LineBuffer2(1457);
--            LineBuffer2(1459) <= LineBuffer2(1458);    
--            LineBuffer2(1460) <= LineBuffer2(1459);
--            LineBuffer2(1461) <= LineBuffer2(1460);
--            LineBuffer2(1462) <= LineBuffer2(1461);
--            LineBuffer2(1463) <= LineBuffer2(1462);
--            LineBuffer2(1464) <= LineBuffer2(1463);
--            LineBuffer2(1465) <= LineBuffer2(1464);
--            LineBuffer2(1466) <= LineBuffer2(1465);
--            LineBuffer2(1467) <= LineBuffer2(1466);
--            LineBuffer2(1468) <= LineBuffer2(1467);
--            LineBuffer2(1469) <= LineBuffer2(1468);    
--            LineBuffer2(1470) <= LineBuffer2(1469);
--            LineBuffer2(1471) <= LineBuffer2(1470);
--            LineBuffer2(1472) <= LineBuffer2(1471);
--            LineBuffer2(1473) <= LineBuffer2(1472);
--            LineBuffer2(1474) <= LineBuffer2(1473);
--            LineBuffer2(1475) <= LineBuffer2(1474);
--            LineBuffer2(1476) <= LineBuffer2(1475);
--            LineBuffer2(1477) <= LineBuffer2(1476);
--            LineBuffer2(1478) <= LineBuffer2(1477);
--            LineBuffer2(1479) <= LineBuffer2(1478);
--            LineBuffer2(1480) <= LineBuffer2(1479);
--            LineBuffer2(1481) <= LineBuffer2(1480);
--            LineBuffer2(1482) <= LineBuffer2(1481);
--            LineBuffer2(1483) <= LineBuffer2(1482);
--            LineBuffer2(1484) <= LineBuffer2(1483);
--            LineBuffer2(1485) <= LineBuffer2(1484);
--            LineBuffer2(1486) <= LineBuffer2(1485);
--            LineBuffer2(1487) <= LineBuffer2(1486);
--            LineBuffer2(1488) <= LineBuffer2(1487);
--            LineBuffer2(1489) <= LineBuffer2(1488);    
--            LineBuffer2(1490) <= LineBuffer2(1489);
--            LineBuffer2(1491) <= LineBuffer2(1490);
--            LineBuffer2(1492) <= LineBuffer2(1491);
--            LineBuffer2(1493) <= LineBuffer2(1492);
--            LineBuffer2(1494) <= LineBuffer2(1493);
--            LineBuffer2(1495) <= LineBuffer2(1494);
--            LineBuffer2(1496) <= LineBuffer2(1495);
--            LineBuffer2(1497) <= LineBuffer2(1496);
--            LineBuffer2(1498) <= LineBuffer2(1497);
--            LineBuffer2(1499) <= LineBuffer2(1498);    
--            LineBuffer2(1500) <= LineBuffer2(1499);
--            LineBuffer2(1501) <= LineBuffer2(1500);
--            LineBuffer2(1502) <= LineBuffer2(1501);
--            LineBuffer2(1503) <= LineBuffer2(1502);
--            LineBuffer2(1504) <= LineBuffer2(1503);
--            LineBuffer2(1505) <= LineBuffer2(1504);
--            LineBuffer2(1506) <= LineBuffer2(1505);
--            LineBuffer2(1507) <= LineBuffer2(1506);
--            LineBuffer2(1508) <= LineBuffer2(1507);
--            LineBuffer2(1509) <= LineBuffer2(1508);    
--            LineBuffer2(1510) <= LineBuffer2(1509);
--            LineBuffer2(1511) <= LineBuffer2(1510);
--            LineBuffer2(1512) <= LineBuffer2(1511);
--            LineBuffer2(1513) <= LineBuffer2(1512);
--            LineBuffer2(1514) <= LineBuffer2(1513);
--            LineBuffer2(1515) <= LineBuffer2(1514);
--            LineBuffer2(1516) <= LineBuffer2(1515);
--            LineBuffer2(1517) <= LineBuffer2(1516);
--            LineBuffer2(1518) <= LineBuffer2(1517);
--            LineBuffer2(1519) <= LineBuffer2(1518);    
--            LineBuffer2(1520) <= LineBuffer2(1519);
--            LineBuffer2(1521) <= LineBuffer2(1520);
--            LineBuffer2(1522) <= LineBuffer2(1521);
--            LineBuffer2(1523) <= LineBuffer2(1522);
--            LineBuffer2(1524) <= LineBuffer2(1523);
--            LineBuffer2(1525) <= LineBuffer2(1524);
--            LineBuffer2(1526) <= LineBuffer2(1525);
--            LineBuffer2(1527) <= LineBuffer2(1526);
--            LineBuffer2(1528) <= LineBuffer2(1527);
--            LineBuffer2(1529) <= LineBuffer2(1528);    
--            LineBuffer2(1530) <= LineBuffer2(1529);
--            LineBuffer2(1531) <= LineBuffer2(1530);
--            LineBuffer2(1532) <= LineBuffer2(1531);
--            LineBuffer2(1533) <= LineBuffer2(1532);
--            LineBuffer2(1534) <= LineBuffer2(1533);
--            LineBuffer2(1535) <= LineBuffer2(1534);
--            LineBuffer2(1536) <= LineBuffer2(1535);
--            LineBuffer2(1537) <= LineBuffer2(1536);
--            LineBuffer2(1538) <= LineBuffer2(1537);
--            LineBuffer2(1539) <= LineBuffer2(1538);    
--            LineBuffer2(1540) <= LineBuffer2(1539);
--            LineBuffer2(1541) <= LineBuffer2(1540);
--            LineBuffer2(1542) <= LineBuffer2(1541);
--            LineBuffer2(1543) <= LineBuffer2(1542);
--            LineBuffer2(1544) <= LineBuffer2(1543);
--            LineBuffer2(1545) <= LineBuffer2(1544);
--            LineBuffer2(1546) <= LineBuffer2(1545);
--            LineBuffer2(1547) <= LineBuffer2(1546);
--            LineBuffer2(1548) <= LineBuffer2(1547);
--            LineBuffer2(1549) <= LineBuffer2(1548);    
--            LineBuffer2(1550) <= LineBuffer2(1549);
--            LineBuffer2(1551) <= LineBuffer2(1550);
--            LineBuffer2(1552) <= LineBuffer2(1551);
--            LineBuffer2(1553) <= LineBuffer2(1552);
--            LineBuffer2(1554) <= LineBuffer2(1553);
--            LineBuffer2(1555) <= LineBuffer2(1554);
--            LineBuffer2(1556) <= LineBuffer2(1555);
--            LineBuffer2(1557) <= LineBuffer2(1556);
--            LineBuffer2(1558) <= LineBuffer2(1557);
--            LineBuffer2(1559) <= LineBuffer2(1558);    
--            LineBuffer2(1560) <= LineBuffer2(1559);
--            LineBuffer2(1561) <= LineBuffer2(1560);
--            LineBuffer2(1562) <= LineBuffer2(1561);
--            LineBuffer2(1563) <= LineBuffer2(1562);
--            LineBuffer2(1564) <= LineBuffer2(1563);
--            LineBuffer2(1565) <= LineBuffer2(1564);
--            LineBuffer2(1566) <= LineBuffer2(1565);
--            LineBuffer2(1567) <= LineBuffer2(1566);
--            LineBuffer2(1568) <= LineBuffer2(1567);
--            LineBuffer2(1569) <= LineBuffer2(1568);    
--            LineBuffer2(1570) <= LineBuffer2(1569);
--            LineBuffer2(1571) <= LineBuffer2(1570);
--            LineBuffer2(1572) <= LineBuffer2(1571);
--            LineBuffer2(1573) <= LineBuffer2(1572);
--            LineBuffer2(1574) <= LineBuffer2(1573);
--            LineBuffer2(1575) <= LineBuffer2(1574);
--            LineBuffer2(1576) <= LineBuffer2(1575);
--            LineBuffer2(1577) <= LineBuffer2(1576);
--            LineBuffer2(1578) <= LineBuffer2(1577);
--            LineBuffer2(1579) <= LineBuffer2(1578);
--            LineBuffer2(1580) <= LineBuffer2(1579);
--            LineBuffer2(1581) <= LineBuffer2(1580);
--            LineBuffer2(1582) <= LineBuffer2(1581);
--            LineBuffer2(1583) <= LineBuffer2(1582);
--            LineBuffer2(1584) <= LineBuffer2(1583);
--            LineBuffer2(1585) <= LineBuffer2(1584);
--            LineBuffer2(1586) <= LineBuffer2(1585);
--            LineBuffer2(1587) <= LineBuffer2(1586);
--            LineBuffer2(1588) <= LineBuffer2(1587);
--            LineBuffer2(1589) <= LineBuffer2(1588);    
--            LineBuffer2(1590) <= LineBuffer2(1589);
--            LineBuffer2(1591) <= LineBuffer2(1590);
--            LineBuffer2(1592) <= LineBuffer2(1591);
--            LineBuffer2(1593) <= LineBuffer2(1592);
--            LineBuffer2(1594) <= LineBuffer2(1593);
--            LineBuffer2(1595) <= LineBuffer2(1594);
--            LineBuffer2(1596) <= LineBuffer2(1595);
--            LineBuffer2(1597) <= LineBuffer2(1596);
--            LineBuffer2(1598) <= LineBuffer2(1597);
--            LineBuffer2(1599) <= LineBuffer2(1598);    
--            LineBuffer2(1600) <= LineBuffer2(1599);
--            LineBuffer2(1601) <= LineBuffer2(1600);
--            LineBuffer2(1602) <= LineBuffer2(1601);
--            LineBuffer2(1603) <= LineBuffer2(1602);
--            LineBuffer2(1604) <= LineBuffer2(1603);
--            LineBuffer2(1605) <= LineBuffer2(1604);
--            LineBuffer2(1606) <= LineBuffer2(1605);
--            LineBuffer2(1607) <= LineBuffer2(1606);
--            LineBuffer2(1608) <= LineBuffer2(1607);
--            LineBuffer2(1609) <= LineBuffer2(1608);    
--            LineBuffer2(1610) <= LineBuffer2(1609);
--            LineBuffer2(1611) <= LineBuffer2(1610);
--            LineBuffer2(1612) <= LineBuffer2(1611);
--            LineBuffer2(1613) <= LineBuffer2(1612);
--            LineBuffer2(1614) <= LineBuffer2(1613);
--            LineBuffer2(1615) <= LineBuffer2(1614);
--            LineBuffer2(1616) <= LineBuffer2(1615);
--            LineBuffer2(1617) <= LineBuffer2(1616);
--            LineBuffer2(1618) <= LineBuffer2(1617);
--            LineBuffer2(1619) <= LineBuffer2(1618);    
--            LineBuffer2(1620) <= LineBuffer2(1619);
--            LineBuffer2(1621) <= LineBuffer2(1620);
--            LineBuffer2(1622) <= LineBuffer2(1621);
--            LineBuffer2(1623) <= LineBuffer2(1622);
--            LineBuffer2(1624) <= LineBuffer2(1623);
--            LineBuffer2(1625) <= LineBuffer2(1624);
--            LineBuffer2(1626) <= LineBuffer2(1625);
--            LineBuffer2(1627) <= LineBuffer2(1626);
--            LineBuffer2(1628) <= LineBuffer2(1627);
--            LineBuffer2(1629) <= LineBuffer2(1628);    
--            LineBuffer2(1630) <= LineBuffer2(1629);
--            LineBuffer2(1631) <= LineBuffer2(1630);
--            LineBuffer2(1632) <= LineBuffer2(1631);
--            LineBuffer2(1633) <= LineBuffer2(1632);
--            LineBuffer2(1634) <= LineBuffer2(1633);
--            LineBuffer2(1635) <= LineBuffer2(1634);
--            LineBuffer2(1636) <= LineBuffer2(1635);
--            LineBuffer2(1637) <= LineBuffer2(1636);
--            LineBuffer2(1638) <= LineBuffer2(1637);
--            LineBuffer2(1639) <= LineBuffer2(1638);    
--            LineBuffer2(1640) <= LineBuffer2(1639);
--            LineBuffer2(1641) <= LineBuffer2(1640);
--            LineBuffer2(1642) <= LineBuffer2(1641);
--            LineBuffer2(1643) <= LineBuffer2(1642);
--            LineBuffer2(1644) <= LineBuffer2(1643);
--            LineBuffer2(1645) <= LineBuffer2(1644);
--            LineBuffer2(1646) <= LineBuffer2(1645);
--            LineBuffer2(1647) <= LineBuffer2(1646);
--            LineBuffer2(1648) <= LineBuffer2(1647);
--            LineBuffer2(1649) <= LineBuffer2(1648);    
--            LineBuffer2(1650) <= LineBuffer2(1649);
--            LineBuffer2(1651) <= LineBuffer2(1650);
--            LineBuffer2(1652) <= LineBuffer2(1651);
--            LineBuffer2(1653) <= LineBuffer2(1652);
--            LineBuffer2(1654) <= LineBuffer2(1653);
--            LineBuffer2(1655) <= LineBuffer2(1654);
--            LineBuffer2(1656) <= LineBuffer2(1655);
--            LineBuffer2(1657) <= LineBuffer2(1656);
--            LineBuffer2(1658) <= LineBuffer2(1657);
--            LineBuffer2(1659) <= LineBuffer2(1658);    
--            LineBuffer2(1660) <= LineBuffer2(1659);
--            LineBuffer2(1661) <= LineBuffer2(1660);
--            LineBuffer2(1662) <= LineBuffer2(1661);
--            LineBuffer2(1663) <= LineBuffer2(1662);
--            LineBuffer2(1664) <= LineBuffer2(1663);
--            LineBuffer2(1665) <= LineBuffer2(1664);
--            LineBuffer2(1666) <= LineBuffer2(1665);
--            LineBuffer2(1667) <= LineBuffer2(1666);
--            LineBuffer2(1668) <= LineBuffer2(1667);
--            LineBuffer2(1669) <= LineBuffer2(1668);    
--            LineBuffer2(1670) <= LineBuffer2(1669);
--            LineBuffer2(1671) <= LineBuffer2(1670);
--            LineBuffer2(1672) <= LineBuffer2(1671);
--            LineBuffer2(1673) <= LineBuffer2(1672);
--            LineBuffer2(1674) <= LineBuffer2(1673);
--            LineBuffer2(1675) <= LineBuffer2(1674);
--            LineBuffer2(1676) <= LineBuffer2(1675);
--            LineBuffer2(1677) <= LineBuffer2(1676);
--            LineBuffer2(1678) <= LineBuffer2(1677);
--            LineBuffer2(1679) <= LineBuffer2(1678);
--            LineBuffer2(1680) <= LineBuffer2(1679);
--            LineBuffer2(1681) <= LineBuffer2(1680);
--            LineBuffer2(1682) <= LineBuffer2(1681);
--            LineBuffer2(1683) <= LineBuffer2(1682);
--            LineBuffer2(1684) <= LineBuffer2(1683);
--            LineBuffer2(1685) <= LineBuffer2(1684);
--            LineBuffer2(1686) <= LineBuffer2(1685);
--            LineBuffer2(1687) <= LineBuffer2(1686);
--            LineBuffer2(1688) <= LineBuffer2(1687);
--            LineBuffer2(1689) <= LineBuffer2(1688);    
--            LineBuffer2(1690) <= LineBuffer2(1689);
--            LineBuffer2(1691) <= LineBuffer2(1690);
--            LineBuffer2(1692) <= LineBuffer2(1691);
--            LineBuffer2(1693) <= LineBuffer2(1692);
--            LineBuffer2(1694) <= LineBuffer2(1693);
--            LineBuffer2(1695) <= LineBuffer2(1694);
--            LineBuffer2(1696) <= LineBuffer2(1695);
--            LineBuffer2(1697) <= LineBuffer2(1696);
--            LineBuffer2(1698) <= LineBuffer2(1697);
--            LineBuffer2(1699) <= LineBuffer2(1698);    
--            LineBuffer2(1700) <= LineBuffer2(1699);
--            LineBuffer2(1701) <= LineBuffer2(1700);
--            LineBuffer2(1702) <= LineBuffer2(1701);
--            LineBuffer2(1703) <= LineBuffer2(1702);
--            LineBuffer2(1704) <= LineBuffer2(1703);
--            LineBuffer2(1705) <= LineBuffer2(1704);
--            LineBuffer2(1706) <= LineBuffer2(1705);
--            LineBuffer2(1707) <= LineBuffer2(1706);
--            LineBuffer2(1708) <= LineBuffer2(1707);
--            LineBuffer2(1709) <= LineBuffer2(1708);    
--            LineBuffer2(1710) <= LineBuffer2(1709);
--            LineBuffer2(1711) <= LineBuffer2(1710);
--            LineBuffer2(1712) <= LineBuffer2(1711);
--            LineBuffer2(1713) <= LineBuffer2(1712);
--            LineBuffer2(1714) <= LineBuffer2(1713);
--            LineBuffer2(1715) <= LineBuffer2(1714);
--            LineBuffer2(1716) <= LineBuffer2(1715);
--            LineBuffer2(1717) <= LineBuffer2(1716);
--            LineBuffer2(1718) <= LineBuffer2(1717);
--            LineBuffer2(1719) <= LineBuffer2(1718);    
--            LineBuffer2(1720) <= LineBuffer2(1719);
--            LineBuffer2(1721) <= LineBuffer2(1720);
--            LineBuffer2(1722) <= LineBuffer2(1721);
--            LineBuffer2(1723) <= LineBuffer2(1722);
--            LineBuffer2(1724) <= LineBuffer2(1723);
--            LineBuffer2(1725) <= LineBuffer2(1724);
--            LineBuffer2(1726) <= LineBuffer2(1725);
--            LineBuffer2(1727) <= LineBuffer2(1726);
--            LineBuffer2(1728) <= LineBuffer2(1727);
--            LineBuffer2(1729) <= LineBuffer2(1728);    
--            LineBuffer2(1730) <= LineBuffer2(1729);
--            LineBuffer2(1731) <= LineBuffer2(1730);
--            LineBuffer2(1732) <= LineBuffer2(1731);
--            LineBuffer2(1733) <= LineBuffer2(1732);
--            LineBuffer2(1734) <= LineBuffer2(1733);
--            LineBuffer2(1735) <= LineBuffer2(1734);
--            LineBuffer2(1736) <= LineBuffer2(1735);
--            LineBuffer2(1737) <= LineBuffer2(1736);
--            LineBuffer2(1738) <= LineBuffer2(1737);
--            LineBuffer2(1739) <= LineBuffer2(1738);    
--            LineBuffer2(1740) <= LineBuffer2(1739);
--            LineBuffer2(1741) <= LineBuffer2(1740);
--            LineBuffer2(1742) <= LineBuffer2(1741);
--            LineBuffer2(1743) <= LineBuffer2(1742);
--            LineBuffer2(1744) <= LineBuffer2(1743);
--            LineBuffer2(1745) <= LineBuffer2(1744);
--            LineBuffer2(1746) <= LineBuffer2(1745);
--            LineBuffer2(1747) <= LineBuffer2(1746);
--            LineBuffer2(1748) <= LineBuffer2(1747);
--            LineBuffer2(1749) <= LineBuffer2(1748);    
--            LineBuffer2(1750) <= LineBuffer2(1749);
--            LineBuffer2(1751) <= LineBuffer2(1750);
--            LineBuffer2(1752) <= LineBuffer2(1751);
--            LineBuffer2(1753) <= LineBuffer2(1752);
--            LineBuffer2(1754) <= LineBuffer2(1753);
--            LineBuffer2(1755) <= LineBuffer2(1754);
--            LineBuffer2(1756) <= LineBuffer2(1755);
--            LineBuffer2(1757) <= LineBuffer2(1756);
--            LineBuffer2(1758) <= LineBuffer2(1757);
--            LineBuffer2(1759) <= LineBuffer2(1758);    
--            LineBuffer2(1760) <= LineBuffer2(1759);
--            LineBuffer2(1761) <= LineBuffer2(1760);
--            LineBuffer2(1762) <= LineBuffer2(1761);
--            LineBuffer2(1763) <= LineBuffer2(1762);
--            LineBuffer2(1764) <= LineBuffer2(1763);
--            LineBuffer2(1765) <= LineBuffer2(1764);
--            LineBuffer2(1766) <= LineBuffer2(1765);
--            LineBuffer2(1767) <= LineBuffer2(1766);
--            LineBuffer2(1768) <= LineBuffer2(1767);
--            LineBuffer2(1769) <= LineBuffer2(1768);    
--            LineBuffer2(1770) <= LineBuffer2(1769);
--            LineBuffer2(1771) <= LineBuffer2(1770);
--            LineBuffer2(1772) <= LineBuffer2(1771);
--            LineBuffer2(1773) <= LineBuffer2(1772);
--            LineBuffer2(1774) <= LineBuffer2(1773);
--            LineBuffer2(1775) <= LineBuffer2(1774);
--            LineBuffer2(1776) <= LineBuffer2(1775);
--            LineBuffer2(1777) <= LineBuffer2(1776);
--            LineBuffer2(1778) <= LineBuffer2(1777);
--            LineBuffer2(1779) <= LineBuffer2(1778);
--            LineBuffer2(1780) <= LineBuffer2(1779);
--            LineBuffer2(1781) <= LineBuffer2(1780);
--            LineBuffer2(1782) <= LineBuffer2(1781);
--            LineBuffer2(1783) <= LineBuffer2(1782);
--            LineBuffer2(1784) <= LineBuffer2(1783);
--            LineBuffer2(1785) <= LineBuffer2(1784);
--            LineBuffer2(1786) <= LineBuffer2(1785);
--            LineBuffer2(1787) <= LineBuffer2(1786);
--            LineBuffer2(1788) <= LineBuffer2(1787);
--            LineBuffer2(1789) <= LineBuffer2(1788);    
--            LineBuffer2(1790) <= LineBuffer2(1789);
--            LineBuffer2(1791) <= LineBuffer2(1790);
--            LineBuffer2(1792) <= LineBuffer2(1791);
--            LineBuffer2(1793) <= LineBuffer2(1792);
--            LineBuffer2(1794) <= LineBuffer2(1793);
--            LineBuffer2(1795) <= LineBuffer2(1794);
--            LineBuffer2(1796) <= LineBuffer2(1795);
--            LineBuffer2(1797) <= LineBuffer2(1796);
--            LineBuffer2(1798) <= LineBuffer2(1797);
--            LineBuffer2(1799) <= LineBuffer2(1798);    
--            LineBuffer2(1800) <= LineBuffer2(1799);
--            LineBuffer2(1801) <= LineBuffer2(1800);
--            LineBuffer2(1802) <= LineBuffer2(1801);
--            LineBuffer2(1803) <= LineBuffer2(1802);
--            LineBuffer2(1804) <= LineBuffer2(1803);
--            LineBuffer2(1805) <= LineBuffer2(1804);
--            LineBuffer2(1806) <= LineBuffer2(1805);
--            LineBuffer2(1807) <= LineBuffer2(1806);
--            LineBuffer2(1808) <= LineBuffer2(1807);
--            LineBuffer2(1809) <= LineBuffer2(1808);    
--            LineBuffer2(1810) <= LineBuffer2(1809);
--            LineBuffer2(1811) <= LineBuffer2(1810);
--            LineBuffer2(1812) <= LineBuffer2(1811);
--            LineBuffer2(1813) <= LineBuffer2(1812);
--            LineBuffer2(1814) <= LineBuffer2(1813);
--            LineBuffer2(1815) <= LineBuffer2(1814);
--            LineBuffer2(1816) <= LineBuffer2(1815);
--            LineBuffer2(1817) <= LineBuffer2(1816);
--            LineBuffer2(1818) <= LineBuffer2(1817);
--            LineBuffer2(1819) <= LineBuffer2(1818);    
--            LineBuffer2(1820) <= LineBuffer2(1819);
--            LineBuffer2(1821) <= LineBuffer2(1820);
--            LineBuffer2(1822) <= LineBuffer2(1821);
--            LineBuffer2(1823) <= LineBuffer2(1822);
--            LineBuffer2(1824) <= LineBuffer2(1823);
--            LineBuffer2(1825) <= LineBuffer2(1824);
--            LineBuffer2(1826) <= LineBuffer2(1825);
--            LineBuffer2(1827) <= LineBuffer2(1826);
--            LineBuffer2(1828) <= LineBuffer2(1827);
--            LineBuffer2(1829) <= LineBuffer2(1828);    
--            LineBuffer2(1830) <= LineBuffer2(1829);
--            LineBuffer2(1831) <= LineBuffer2(1830);
--            LineBuffer2(1832) <= LineBuffer2(1831);
--            LineBuffer2(1833) <= LineBuffer2(1832);
--            LineBuffer2(1834) <= LineBuffer2(1833);
--            LineBuffer2(1835) <= LineBuffer2(1834);
--            LineBuffer2(1836) <= LineBuffer2(1835);
--            LineBuffer2(1837) <= LineBuffer2(1836);
--            LineBuffer2(1838) <= LineBuffer2(1837);
--            LineBuffer2(1839) <= LineBuffer2(1838);    
--            LineBuffer2(1840) <= LineBuffer2(1839);
--            LineBuffer2(1841) <= LineBuffer2(1840);
--            LineBuffer2(1842) <= LineBuffer2(1841);
--            LineBuffer2(1843) <= LineBuffer2(1842);
--            LineBuffer2(1844) <= LineBuffer2(1843);
--            LineBuffer2(1845) <= LineBuffer2(1844);
--            LineBuffer2(1846) <= LineBuffer2(1845);
--            LineBuffer2(1847) <= LineBuffer2(1846);
--            LineBuffer2(1848) <= LineBuffer2(1847);
--            LineBuffer2(1849) <= LineBuffer2(1848);    
--            LineBuffer2(1850) <= LineBuffer2(1849);
--            LineBuffer2(1851) <= LineBuffer2(1850);
--            LineBuffer2(1852) <= LineBuffer2(1851);
--            LineBuffer2(1853) <= LineBuffer2(1852);
--            LineBuffer2(1854) <= LineBuffer2(1853);
--            LineBuffer2(1855) <= LineBuffer2(1854);
--            LineBuffer2(1856) <= LineBuffer2(1855);
--            LineBuffer2(1857) <= LineBuffer2(1856);
--            LineBuffer2(1858) <= LineBuffer2(1857);
--            LineBuffer2(1859) <= LineBuffer2(1858);    
--            LineBuffer2(1860) <= LineBuffer2(1859);
--            LineBuffer2(1861) <= LineBuffer2(1860);
--            LineBuffer2(1862) <= LineBuffer2(1861);
--            LineBuffer2(1863) <= LineBuffer2(1862);
--            LineBuffer2(1864) <= LineBuffer2(1863);
--            LineBuffer2(1865) <= LineBuffer2(1864);
--            LineBuffer2(1866) <= LineBuffer2(1865);
--            LineBuffer2(1867) <= LineBuffer2(1866);
--            LineBuffer2(1868) <= LineBuffer2(1867);
--            LineBuffer2(1869) <= LineBuffer2(1868);    
--            LineBuffer2(1870) <= LineBuffer2(1869);
--            LineBuffer2(1871) <= LineBuffer2(1870);
--            LineBuffer2(1872) <= LineBuffer2(1871);
--            LineBuffer2(1873) <= LineBuffer2(1872);
--            LineBuffer2(1874) <= LineBuffer2(1873);
--            LineBuffer2(1875) <= LineBuffer2(1874);
--            LineBuffer2(1876) <= LineBuffer2(1875);
--            LineBuffer2(1877) <= LineBuffer2(1876);
--            LineBuffer2(1878) <= LineBuffer2(1877);
--            LineBuffer2(1879) <= LineBuffer2(1878);
--            LineBuffer2(1880) <= LineBuffer2(1879);
--            LineBuffer2(1881) <= LineBuffer2(1880);
--            LineBuffer2(1882) <= LineBuffer2(1881);
--            LineBuffer2(1883) <= LineBuffer2(1882);
--            LineBuffer2(1884) <= LineBuffer2(1883);
--            LineBuffer2(1885) <= LineBuffer2(1884);
--            LineBuffer2(1886) <= LineBuffer2(1885);
--            LineBuffer2(1887) <= LineBuffer2(1886);
--            LineBuffer2(1888) <= LineBuffer2(1887);
--            LineBuffer2(1889) <= LineBuffer2(1888);    
--            LineBuffer2(1890) <= LineBuffer2(1889);
--            LineBuffer2(1891) <= LineBuffer2(1890);
--            LineBuffer2(1892) <= LineBuffer2(1891);
--            LineBuffer2(1893) <= LineBuffer2(1892);
--            LineBuffer2(1894) <= LineBuffer2(1893);
--            LineBuffer2(1895) <= LineBuffer2(1894);
--            LineBuffer2(1896) <= LineBuffer2(1895);
--            LineBuffer2(1897) <= LineBuffer2(1896);
--            LineBuffer2(1898) <= LineBuffer2(1897);
--            LineBuffer2(1899) <= LineBuffer2(1898);    
--            LineBuffer2(1900) <= LineBuffer2(1899);
--            LineBuffer2(1901) <= LineBuffer2(1900);
--            LineBuffer2(1902) <= LineBuffer2(1901);
--            LineBuffer2(1903) <= LineBuffer2(1902);
--            LineBuffer2(1904) <= LineBuffer2(1903);
--            LineBuffer2(1905) <= LineBuffer2(1904);
--            LineBuffer2(1906) <= LineBuffer2(1905);
--            LineBuffer2(1907) <= LineBuffer2(1906);
--            LineBuffer2(1908) <= LineBuffer2(1907);
--            LineBuffer2(1909) <= LineBuffer2(1908);    
--            LineBuffer2(1910) <= LineBuffer2(1909);
--            LineBuffer2(1911) <= LineBuffer2(1910);
--            LineBuffer2(1912) <= LineBuffer2(1911);
--            LineBuffer2(1913) <= LineBuffer2(1912);
--            LineBuffer2(1914) <= LineBuffer2(1913);
--            LineBuffer2(1915) <= LineBuffer2(1914);
--            LineBuffer2(1916) <= LineBuffer2(1915);
--            LineBuffer2(1917) <= LineBuffer2(1916);
--            LineBuffer2(1918) <= LineBuffer2(1917);
--            LineBuffer2(1919) <= LineBuffer2(1918);					
			end if;
	end if;
 end if;
end process;

taps_signal(23 downto 0) <= LineBuffer2(1279) & LineBuffer1(1279) & LineBuffer0(1279);
shiftout(7 downto 0) <= LineBuffer2(1279);
taps(23 downto 0) <= taps_signal(23 downto 0);
end Behavioral;
